magic
tech sky130A
magscale 1 2
timestamp 1623636542
<< nwell >>
rect 562120 494182 567614 495550
rect 502426 460824 505768 470352
rect 503026 454632 510928 460552
rect 503028 453842 510928 454632
rect 562120 453880 567614 455248
rect 503026 449132 510928 453842
rect 503028 448342 510928 449132
rect 503026 443174 510928 448342
rect 503026 442286 510926 443174
<< pwell >>
rect 572280 494226 577774 495584
rect 572280 453924 577774 455282
rect 503344 438355 513700 438508
rect 503344 437321 503497 438355
rect 504531 437321 504785 438355
rect 505819 437321 506073 438355
rect 507107 437321 507361 438355
rect 508395 437321 508649 438355
rect 509683 437321 509937 438355
rect 510971 437321 511225 438355
rect 512259 437321 512513 438355
rect 513547 437321 513700 438355
rect 503344 437067 513700 437321
rect 503344 436033 503497 437067
rect 504531 436033 504785 437067
rect 505819 436033 506073 437067
rect 507107 436033 507361 437067
rect 508395 436033 508649 437067
rect 509683 436033 509937 437067
rect 510971 436033 511225 437067
rect 512259 436033 512513 437067
rect 513547 436033 513700 437067
rect 503344 435779 513700 436033
rect 503344 434745 503497 435779
rect 504531 434745 504785 435779
rect 505819 434745 506073 435779
rect 507107 434745 507361 435779
rect 508395 434745 508649 435779
rect 509683 434745 509937 435779
rect 510971 434745 511225 435779
rect 512259 434745 512513 435779
rect 513547 434745 513700 435779
rect 503344 434491 513700 434745
rect 503344 433457 503497 434491
rect 504531 433457 504785 434491
rect 505819 433457 506073 434491
rect 507107 433457 507361 434491
rect 508395 433457 508649 434491
rect 509683 433457 509937 434491
rect 510971 433457 511225 434491
rect 512259 433457 512513 434491
rect 513547 433457 513700 434491
rect 503344 433203 513700 433457
rect 503344 432169 503497 433203
rect 504531 432169 504785 433203
rect 505819 432169 506073 433203
rect 507107 432169 507361 433203
rect 508395 432169 508649 433203
rect 509683 432169 509937 433203
rect 510971 432169 511225 433203
rect 512259 432169 512513 433203
rect 513547 432169 513700 433203
rect 503344 432016 513700 432169
<< nbase >>
rect 503497 437321 504531 438355
rect 504785 437321 505819 438355
rect 506073 437321 507107 438355
rect 507361 437321 508395 438355
rect 508649 437321 509683 438355
rect 509937 437321 510971 438355
rect 511225 437321 512259 438355
rect 512513 437321 513547 438355
rect 503497 436033 504531 437067
rect 504785 436033 505819 437067
rect 506073 436033 507107 437067
rect 507361 436033 508395 437067
rect 508649 436033 509683 437067
rect 509937 436033 510971 437067
rect 511225 436033 512259 437067
rect 512513 436033 513547 437067
rect 503497 434745 504531 435779
rect 504785 434745 505819 435779
rect 506073 434745 507107 435779
rect 507361 434745 508395 435779
rect 508649 434745 509683 435779
rect 509937 434745 510971 435779
rect 511225 434745 512259 435779
rect 512513 434745 513547 435779
rect 503497 433457 504531 434491
rect 504785 433457 505819 434491
rect 506073 433457 507107 434491
rect 507361 433457 508395 434491
rect 508649 433457 509683 434491
rect 509937 433457 510971 434491
rect 511225 433457 512259 434491
rect 512513 433457 513547 434491
rect 503497 432169 504531 433203
rect 504785 432169 505819 433203
rect 506073 432169 507107 433203
rect 507361 432169 508395 433203
rect 508649 432169 509683 433203
rect 509937 432169 510971 433203
rect 511225 432169 512259 433203
rect 512513 432169 513547 433203
<< pmoslvt >>
rect 562316 494402 562516 495402
rect 562574 494402 562774 495402
rect 562832 494402 563032 495402
rect 563090 494402 563290 495402
rect 563348 494402 563548 495402
rect 563606 494402 563806 495402
rect 563864 494402 564064 495402
rect 564122 494402 564322 495402
rect 564380 494402 564580 495402
rect 564638 494402 564838 495402
rect 564896 494402 565096 495402
rect 565154 494402 565354 495402
rect 565412 494402 565612 495402
rect 565670 494402 565870 495402
rect 565928 494402 566128 495402
rect 566186 494402 566386 495402
rect 566444 494402 566644 495402
rect 566702 494402 566902 495402
rect 566960 494402 567160 495402
rect 567218 494402 567418 495402
rect 503088 469114 505668 469514
rect 503088 468542 505668 468942
rect 503088 467970 505668 468370
rect 503088 467398 505668 467798
rect 503088 466826 505668 467226
rect 503088 466254 505668 466654
rect 503088 465682 505668 466082
rect 503088 465110 505668 465510
rect 503088 464538 505668 464938
rect 503088 463966 505668 464366
rect 503088 463394 505668 463794
rect 503088 462822 505668 463222
rect 503088 462250 505668 462650
rect 503088 461678 505668 462078
rect 503126 459306 510866 459706
rect 503126 458848 510866 459248
rect 503126 458390 510866 458790
rect 503126 457932 510866 458332
rect 503126 457474 510866 457874
rect 503126 457016 510866 457416
rect 503126 456558 510866 456958
rect 503126 456100 510866 456500
rect 503126 455642 510866 456042
rect 503126 455184 510866 455584
rect 503126 454726 510866 455126
rect 503126 453348 510866 453748
rect 503126 452890 510866 453290
rect 503126 452432 510866 452832
rect 503126 451974 510866 452374
rect 503126 451516 510866 451916
rect 503126 451058 510866 451458
rect 503126 450600 510866 451000
rect 503126 450142 510866 450542
rect 503126 449684 510866 450084
rect 503126 449226 510866 449626
rect 503126 447848 510866 448248
rect 503126 447390 510866 447790
rect 503126 446932 510866 447332
rect 503126 446474 510866 446874
rect 503126 446016 510866 446416
rect 503126 445558 510866 445958
rect 503126 445100 510866 445500
rect 503126 444642 510866 445042
rect 503126 444184 510866 444584
rect 503126 443726 510866 444126
rect 503126 443268 510866 443668
rect 562316 454100 562516 455100
rect 562574 454100 562774 455100
rect 562832 454100 563032 455100
rect 563090 454100 563290 455100
rect 563348 454100 563548 455100
rect 563606 454100 563806 455100
rect 563864 454100 564064 455100
rect 564122 454100 564322 455100
rect 564380 454100 564580 455100
rect 564638 454100 564838 455100
rect 564896 454100 565096 455100
rect 565154 454100 565354 455100
rect 565412 454100 565612 455100
rect 565670 454100 565870 455100
rect 565928 454100 566128 455100
rect 566186 454100 566386 455100
rect 566444 454100 566644 455100
rect 566702 454100 566902 455100
rect 566960 454100 567160 455100
rect 567218 454100 567418 455100
<< nmoslvt >>
rect 572476 494436 572676 495436
rect 572734 494436 572934 495436
rect 572992 494436 573192 495436
rect 573250 494436 573450 495436
rect 573508 494436 573708 495436
rect 573766 494436 573966 495436
rect 574024 494436 574224 495436
rect 574282 494436 574482 495436
rect 574540 494436 574740 495436
rect 574798 494436 574998 495436
rect 575056 494436 575256 495436
rect 575314 494436 575514 495436
rect 575572 494436 575772 495436
rect 575830 494436 576030 495436
rect 576088 494436 576288 495436
rect 576346 494436 576546 495436
rect 576604 494436 576804 495436
rect 576862 494436 577062 495436
rect 577120 494436 577320 495436
rect 577378 494436 577578 495436
rect 506558 472318 506958 472718
rect 506558 471860 506958 472260
rect 506558 471402 506958 471802
rect 506558 470944 506958 471344
rect 506558 470486 506958 470886
rect 506558 470028 506958 470428
rect 506280 467388 508080 467788
rect 506280 466816 508080 467216
rect 506280 466244 508080 466644
rect 506280 465672 508080 466072
rect 506280 465100 508080 465500
rect 506280 464528 508080 464928
rect 506280 463956 508080 464356
rect 506280 463384 508080 463784
rect 509832 462728 510232 468128
rect 572476 454134 572676 455134
rect 572734 454134 572934 455134
rect 572992 454134 573192 455134
rect 573250 454134 573450 455134
rect 573508 454134 573708 455134
rect 573766 454134 573966 455134
rect 574024 454134 574224 455134
rect 574282 454134 574482 455134
rect 574540 454134 574740 455134
rect 574798 454134 574998 455134
rect 575056 454134 575256 455134
rect 575314 454134 575514 455134
rect 575572 454134 575772 455134
rect 575830 454134 576030 455134
rect 576088 454134 576288 455134
rect 576346 454134 576546 455134
rect 576604 454134 576804 455134
rect 576862 454134 577062 455134
rect 577120 454134 577320 455134
rect 577378 454134 577578 455134
<< ndiff >>
rect 572418 495424 572476 495436
rect 572418 494448 572430 495424
rect 572464 494448 572476 495424
rect 572418 494436 572476 494448
rect 572676 495424 572734 495436
rect 572676 494448 572688 495424
rect 572722 494448 572734 495424
rect 572676 494436 572734 494448
rect 572934 495424 572992 495436
rect 572934 494448 572946 495424
rect 572980 494448 572992 495424
rect 572934 494436 572992 494448
rect 573192 495424 573250 495436
rect 573192 494448 573204 495424
rect 573238 494448 573250 495424
rect 573192 494436 573250 494448
rect 573450 495424 573508 495436
rect 573450 494448 573462 495424
rect 573496 494448 573508 495424
rect 573450 494436 573508 494448
rect 573708 495424 573766 495436
rect 573708 494448 573720 495424
rect 573754 494448 573766 495424
rect 573708 494436 573766 494448
rect 573966 495424 574024 495436
rect 573966 494448 573978 495424
rect 574012 494448 574024 495424
rect 573966 494436 574024 494448
rect 574224 495424 574282 495436
rect 574224 494448 574236 495424
rect 574270 494448 574282 495424
rect 574224 494436 574282 494448
rect 574482 495424 574540 495436
rect 574482 494448 574494 495424
rect 574528 494448 574540 495424
rect 574482 494436 574540 494448
rect 574740 495424 574798 495436
rect 574740 494448 574752 495424
rect 574786 494448 574798 495424
rect 574740 494436 574798 494448
rect 574998 495424 575056 495436
rect 574998 494448 575010 495424
rect 575044 494448 575056 495424
rect 574998 494436 575056 494448
rect 575256 495424 575314 495436
rect 575256 494448 575268 495424
rect 575302 494448 575314 495424
rect 575256 494436 575314 494448
rect 575514 495424 575572 495436
rect 575514 494448 575526 495424
rect 575560 494448 575572 495424
rect 575514 494436 575572 494448
rect 575772 495424 575830 495436
rect 575772 494448 575784 495424
rect 575818 494448 575830 495424
rect 575772 494436 575830 494448
rect 576030 495424 576088 495436
rect 576030 494448 576042 495424
rect 576076 494448 576088 495424
rect 576030 494436 576088 494448
rect 576288 495424 576346 495436
rect 576288 494448 576300 495424
rect 576334 494448 576346 495424
rect 576288 494436 576346 494448
rect 576546 495424 576604 495436
rect 576546 494448 576558 495424
rect 576592 494448 576604 495424
rect 576546 494436 576604 494448
rect 576804 495424 576862 495436
rect 576804 494448 576816 495424
rect 576850 494448 576862 495424
rect 576804 494436 576862 494448
rect 577062 495424 577120 495436
rect 577062 494448 577074 495424
rect 577108 494448 577120 495424
rect 577062 494436 577120 494448
rect 577320 495424 577378 495436
rect 577320 494448 577332 495424
rect 577366 494448 577378 495424
rect 577320 494436 577378 494448
rect 577578 495424 577636 495436
rect 577578 494448 577590 495424
rect 577624 494448 577636 495424
rect 577578 494436 577636 494448
rect 506558 472764 506958 472776
rect 506558 472730 506570 472764
rect 506946 472730 506958 472764
rect 506558 472718 506958 472730
rect 506558 472306 506958 472318
rect 506558 472272 506570 472306
rect 506946 472272 506958 472306
rect 506558 472260 506958 472272
rect 506558 471848 506958 471860
rect 506558 471814 506570 471848
rect 506946 471814 506958 471848
rect 506558 471802 506958 471814
rect 506558 471390 506958 471402
rect 506558 471356 506570 471390
rect 506946 471356 506958 471390
rect 506558 471344 506958 471356
rect 506558 470932 506958 470944
rect 506558 470898 506570 470932
rect 506946 470898 506958 470932
rect 506558 470886 506958 470898
rect 506558 470474 506958 470486
rect 506558 470440 506570 470474
rect 506946 470440 506958 470474
rect 506558 470428 506958 470440
rect 506558 470016 506958 470028
rect 506558 469982 506570 470016
rect 506946 469982 506958 470016
rect 506558 469970 506958 469982
rect 509774 468116 509832 468128
rect 506280 467834 508080 467846
rect 506280 467800 506292 467834
rect 508068 467800 508080 467834
rect 506280 467788 508080 467800
rect 506280 467376 508080 467388
rect 506280 467342 506292 467376
rect 508068 467342 508080 467376
rect 506280 467330 508080 467342
rect 506280 467262 508080 467274
rect 506280 467228 506292 467262
rect 508068 467228 508080 467262
rect 506280 467216 508080 467228
rect 506280 466804 508080 466816
rect 506280 466770 506292 466804
rect 508068 466770 508080 466804
rect 506280 466758 508080 466770
rect 506280 466690 508080 466702
rect 506280 466656 506292 466690
rect 508068 466656 508080 466690
rect 506280 466644 508080 466656
rect 506280 466232 508080 466244
rect 506280 466198 506292 466232
rect 508068 466198 508080 466232
rect 506280 466186 508080 466198
rect 506280 466118 508080 466130
rect 506280 466084 506292 466118
rect 508068 466084 508080 466118
rect 506280 466072 508080 466084
rect 506280 465660 508080 465672
rect 506280 465626 506292 465660
rect 508068 465626 508080 465660
rect 506280 465614 508080 465626
rect 506280 465546 508080 465558
rect 506280 465512 506292 465546
rect 508068 465512 508080 465546
rect 506280 465500 508080 465512
rect 506280 465088 508080 465100
rect 506280 465054 506292 465088
rect 508068 465054 508080 465088
rect 506280 465042 508080 465054
rect 506280 464974 508080 464986
rect 506280 464940 506292 464974
rect 508068 464940 508080 464974
rect 506280 464928 508080 464940
rect 506280 464516 508080 464528
rect 506280 464482 506292 464516
rect 508068 464482 508080 464516
rect 506280 464470 508080 464482
rect 506280 464402 508080 464414
rect 506280 464368 506292 464402
rect 508068 464368 508080 464402
rect 506280 464356 508080 464368
rect 506280 463944 508080 463956
rect 506280 463910 506292 463944
rect 508068 463910 508080 463944
rect 506280 463898 508080 463910
rect 506280 463830 508080 463842
rect 506280 463796 506292 463830
rect 508068 463796 508080 463830
rect 506280 463784 508080 463796
rect 506280 463372 508080 463384
rect 506280 463338 506292 463372
rect 508068 463338 508080 463372
rect 506280 463326 508080 463338
rect 509774 462740 509786 468116
rect 509820 462740 509832 468116
rect 509774 462728 509832 462740
rect 510232 468116 510290 468128
rect 510232 462740 510244 468116
rect 510278 462740 510290 468116
rect 510232 462728 510290 462740
rect 572418 455122 572476 455134
rect 572418 454146 572430 455122
rect 572464 454146 572476 455122
rect 572418 454134 572476 454146
rect 572676 455122 572734 455134
rect 572676 454146 572688 455122
rect 572722 454146 572734 455122
rect 572676 454134 572734 454146
rect 572934 455122 572992 455134
rect 572934 454146 572946 455122
rect 572980 454146 572992 455122
rect 572934 454134 572992 454146
rect 573192 455122 573250 455134
rect 573192 454146 573204 455122
rect 573238 454146 573250 455122
rect 573192 454134 573250 454146
rect 573450 455122 573508 455134
rect 573450 454146 573462 455122
rect 573496 454146 573508 455122
rect 573450 454134 573508 454146
rect 573708 455122 573766 455134
rect 573708 454146 573720 455122
rect 573754 454146 573766 455122
rect 573708 454134 573766 454146
rect 573966 455122 574024 455134
rect 573966 454146 573978 455122
rect 574012 454146 574024 455122
rect 573966 454134 574024 454146
rect 574224 455122 574282 455134
rect 574224 454146 574236 455122
rect 574270 454146 574282 455122
rect 574224 454134 574282 454146
rect 574482 455122 574540 455134
rect 574482 454146 574494 455122
rect 574528 454146 574540 455122
rect 574482 454134 574540 454146
rect 574740 455122 574798 455134
rect 574740 454146 574752 455122
rect 574786 454146 574798 455122
rect 574740 454134 574798 454146
rect 574998 455122 575056 455134
rect 574998 454146 575010 455122
rect 575044 454146 575056 455122
rect 574998 454134 575056 454146
rect 575256 455122 575314 455134
rect 575256 454146 575268 455122
rect 575302 454146 575314 455122
rect 575256 454134 575314 454146
rect 575514 455122 575572 455134
rect 575514 454146 575526 455122
rect 575560 454146 575572 455122
rect 575514 454134 575572 454146
rect 575772 455122 575830 455134
rect 575772 454146 575784 455122
rect 575818 454146 575830 455122
rect 575772 454134 575830 454146
rect 576030 455122 576088 455134
rect 576030 454146 576042 455122
rect 576076 454146 576088 455122
rect 576030 454134 576088 454146
rect 576288 455122 576346 455134
rect 576288 454146 576300 455122
rect 576334 454146 576346 455122
rect 576288 454134 576346 454146
rect 576546 455122 576604 455134
rect 576546 454146 576558 455122
rect 576592 454146 576604 455122
rect 576546 454134 576604 454146
rect 576804 455122 576862 455134
rect 576804 454146 576816 455122
rect 576850 454146 576862 455122
rect 576804 454134 576862 454146
rect 577062 455122 577120 455134
rect 577062 454146 577074 455122
rect 577108 454146 577120 455122
rect 577062 454134 577120 454146
rect 577320 455122 577378 455134
rect 577320 454146 577332 455122
rect 577366 454146 577378 455122
rect 577320 454134 577378 454146
rect 577578 455122 577636 455134
rect 577578 454146 577590 455122
rect 577624 454146 577636 455122
rect 577578 454134 577636 454146
<< pdiff >>
rect 562258 495390 562316 495402
rect 562258 494414 562270 495390
rect 562304 494414 562316 495390
rect 562258 494402 562316 494414
rect 562516 495390 562574 495402
rect 562516 494414 562528 495390
rect 562562 494414 562574 495390
rect 562516 494402 562574 494414
rect 562774 495390 562832 495402
rect 562774 494414 562786 495390
rect 562820 494414 562832 495390
rect 562774 494402 562832 494414
rect 563032 495390 563090 495402
rect 563032 494414 563044 495390
rect 563078 494414 563090 495390
rect 563032 494402 563090 494414
rect 563290 495390 563348 495402
rect 563290 494414 563302 495390
rect 563336 494414 563348 495390
rect 563290 494402 563348 494414
rect 563548 495390 563606 495402
rect 563548 494414 563560 495390
rect 563594 494414 563606 495390
rect 563548 494402 563606 494414
rect 563806 495390 563864 495402
rect 563806 494414 563818 495390
rect 563852 494414 563864 495390
rect 563806 494402 563864 494414
rect 564064 495390 564122 495402
rect 564064 494414 564076 495390
rect 564110 494414 564122 495390
rect 564064 494402 564122 494414
rect 564322 495390 564380 495402
rect 564322 494414 564334 495390
rect 564368 494414 564380 495390
rect 564322 494402 564380 494414
rect 564580 495390 564638 495402
rect 564580 494414 564592 495390
rect 564626 494414 564638 495390
rect 564580 494402 564638 494414
rect 564838 495390 564896 495402
rect 564838 494414 564850 495390
rect 564884 494414 564896 495390
rect 564838 494402 564896 494414
rect 565096 495390 565154 495402
rect 565096 494414 565108 495390
rect 565142 494414 565154 495390
rect 565096 494402 565154 494414
rect 565354 495390 565412 495402
rect 565354 494414 565366 495390
rect 565400 494414 565412 495390
rect 565354 494402 565412 494414
rect 565612 495390 565670 495402
rect 565612 494414 565624 495390
rect 565658 494414 565670 495390
rect 565612 494402 565670 494414
rect 565870 495390 565928 495402
rect 565870 494414 565882 495390
rect 565916 494414 565928 495390
rect 565870 494402 565928 494414
rect 566128 495390 566186 495402
rect 566128 494414 566140 495390
rect 566174 494414 566186 495390
rect 566128 494402 566186 494414
rect 566386 495390 566444 495402
rect 566386 494414 566398 495390
rect 566432 494414 566444 495390
rect 566386 494402 566444 494414
rect 566644 495390 566702 495402
rect 566644 494414 566656 495390
rect 566690 494414 566702 495390
rect 566644 494402 566702 494414
rect 566902 495390 566960 495402
rect 566902 494414 566914 495390
rect 566948 494414 566960 495390
rect 566902 494402 566960 494414
rect 567160 495390 567218 495402
rect 567160 494414 567172 495390
rect 567206 494414 567218 495390
rect 567160 494402 567218 494414
rect 567418 495390 567476 495402
rect 567418 494414 567430 495390
rect 567464 494414 567476 495390
rect 567418 494402 567476 494414
rect 503088 469560 505668 469572
rect 503088 469526 503100 469560
rect 505656 469526 505668 469560
rect 503088 469514 505668 469526
rect 503088 469102 505668 469114
rect 503088 469068 503100 469102
rect 505656 469068 505668 469102
rect 503088 469056 505668 469068
rect 503088 468988 505668 469000
rect 503088 468954 503100 468988
rect 505656 468954 505668 468988
rect 503088 468942 505668 468954
rect 503088 468530 505668 468542
rect 503088 468496 503100 468530
rect 505656 468496 505668 468530
rect 503088 468484 505668 468496
rect 503088 468416 505668 468428
rect 503088 468382 503100 468416
rect 505656 468382 505668 468416
rect 503088 468370 505668 468382
rect 503088 467958 505668 467970
rect 503088 467924 503100 467958
rect 505656 467924 505668 467958
rect 503088 467912 505668 467924
rect 503088 467844 505668 467856
rect 503088 467810 503100 467844
rect 505656 467810 505668 467844
rect 503088 467798 505668 467810
rect 503088 467386 505668 467398
rect 503088 467352 503100 467386
rect 505656 467352 505668 467386
rect 503088 467340 505668 467352
rect 503088 467272 505668 467284
rect 503088 467238 503100 467272
rect 505656 467238 505668 467272
rect 503088 467226 505668 467238
rect 503088 466814 505668 466826
rect 503088 466780 503100 466814
rect 505656 466780 505668 466814
rect 503088 466768 505668 466780
rect 503088 466700 505668 466712
rect 503088 466666 503100 466700
rect 505656 466666 505668 466700
rect 503088 466654 505668 466666
rect 503088 466242 505668 466254
rect 503088 466208 503100 466242
rect 505656 466208 505668 466242
rect 503088 466196 505668 466208
rect 503088 466128 505668 466140
rect 503088 466094 503100 466128
rect 505656 466094 505668 466128
rect 503088 466082 505668 466094
rect 503088 465670 505668 465682
rect 503088 465636 503100 465670
rect 505656 465636 505668 465670
rect 503088 465624 505668 465636
rect 503088 465556 505668 465568
rect 503088 465522 503100 465556
rect 505656 465522 505668 465556
rect 503088 465510 505668 465522
rect 503088 465098 505668 465110
rect 503088 465064 503100 465098
rect 505656 465064 505668 465098
rect 503088 465052 505668 465064
rect 503088 464984 505668 464996
rect 503088 464950 503100 464984
rect 505656 464950 505668 464984
rect 503088 464938 505668 464950
rect 503088 464526 505668 464538
rect 503088 464492 503100 464526
rect 505656 464492 505668 464526
rect 503088 464480 505668 464492
rect 503088 464412 505668 464424
rect 503088 464378 503100 464412
rect 505656 464378 505668 464412
rect 503088 464366 505668 464378
rect 503088 463954 505668 463966
rect 503088 463920 503100 463954
rect 505656 463920 505668 463954
rect 503088 463908 505668 463920
rect 503088 463840 505668 463852
rect 503088 463806 503100 463840
rect 505656 463806 505668 463840
rect 503088 463794 505668 463806
rect 503088 463382 505668 463394
rect 503088 463348 503100 463382
rect 505656 463348 505668 463382
rect 503088 463336 505668 463348
rect 503088 463268 505668 463280
rect 503088 463234 503100 463268
rect 505656 463234 505668 463268
rect 503088 463222 505668 463234
rect 503088 462810 505668 462822
rect 503088 462776 503100 462810
rect 505656 462776 505668 462810
rect 503088 462764 505668 462776
rect 503088 462696 505668 462708
rect 503088 462662 503100 462696
rect 505656 462662 505668 462696
rect 503088 462650 505668 462662
rect 503088 462238 505668 462250
rect 503088 462204 503100 462238
rect 505656 462204 505668 462238
rect 503088 462192 505668 462204
rect 503088 462124 505668 462136
rect 503088 462090 503100 462124
rect 505656 462090 505668 462124
rect 503088 462078 505668 462090
rect 503088 461666 505668 461678
rect 503088 461632 503100 461666
rect 505656 461632 505668 461666
rect 503088 461620 505668 461632
rect 503126 459752 510866 459764
rect 503126 459718 503138 459752
rect 510854 459718 510866 459752
rect 503126 459706 510866 459718
rect 503126 459294 510866 459306
rect 503126 459260 503138 459294
rect 510854 459260 510866 459294
rect 503126 459248 510866 459260
rect 503126 458836 510866 458848
rect 503126 458802 503138 458836
rect 510854 458802 510866 458836
rect 503126 458790 510866 458802
rect 503126 458378 510866 458390
rect 503126 458344 503138 458378
rect 510854 458344 510866 458378
rect 503126 458332 510866 458344
rect 503126 457920 510866 457932
rect 503126 457886 503138 457920
rect 510854 457886 510866 457920
rect 503126 457874 510866 457886
rect 503126 457462 510866 457474
rect 503126 457428 503138 457462
rect 510854 457428 510866 457462
rect 503126 457416 510866 457428
rect 503126 457004 510866 457016
rect 503126 456970 503138 457004
rect 510854 456970 510866 457004
rect 503126 456958 510866 456970
rect 503126 456546 510866 456558
rect 503126 456512 503138 456546
rect 510854 456512 510866 456546
rect 503126 456500 510866 456512
rect 503126 456088 510866 456100
rect 503126 456054 503138 456088
rect 510854 456054 510866 456088
rect 503126 456042 510866 456054
rect 503126 455630 510866 455642
rect 503126 455596 503138 455630
rect 510854 455596 510866 455630
rect 503126 455584 510866 455596
rect 503126 455172 510866 455184
rect 503126 455138 503138 455172
rect 510854 455138 510866 455172
rect 503126 455126 510866 455138
rect 503126 454714 510866 454726
rect 503126 454680 503138 454714
rect 510854 454680 510866 454714
rect 503126 454668 510866 454680
rect 503126 453794 510866 453806
rect 503126 453760 503138 453794
rect 510854 453760 510866 453794
rect 503126 453748 510866 453760
rect 503126 453336 510866 453348
rect 503126 453302 503138 453336
rect 510854 453302 510866 453336
rect 503126 453290 510866 453302
rect 503126 452878 510866 452890
rect 503126 452844 503138 452878
rect 510854 452844 510866 452878
rect 503126 452832 510866 452844
rect 503126 452420 510866 452432
rect 503126 452386 503138 452420
rect 510854 452386 510866 452420
rect 503126 452374 510866 452386
rect 503126 451962 510866 451974
rect 503126 451928 503138 451962
rect 510854 451928 510866 451962
rect 503126 451916 510866 451928
rect 503126 451504 510866 451516
rect 503126 451470 503138 451504
rect 510854 451470 510866 451504
rect 503126 451458 510866 451470
rect 503126 451046 510866 451058
rect 503126 451012 503138 451046
rect 510854 451012 510866 451046
rect 503126 451000 510866 451012
rect 503126 450588 510866 450600
rect 503126 450554 503138 450588
rect 510854 450554 510866 450588
rect 503126 450542 510866 450554
rect 503126 450130 510866 450142
rect 503126 450096 503138 450130
rect 510854 450096 510866 450130
rect 503126 450084 510866 450096
rect 503126 449672 510866 449684
rect 503126 449638 503138 449672
rect 510854 449638 510866 449672
rect 503126 449626 510866 449638
rect 503126 449214 510866 449226
rect 503126 449180 503138 449214
rect 510854 449180 510866 449214
rect 503126 449168 510866 449180
rect 503126 448294 510866 448306
rect 503126 448260 503138 448294
rect 510854 448260 510866 448294
rect 503126 448248 510866 448260
rect 503126 447836 510866 447848
rect 503126 447802 503138 447836
rect 510854 447802 510866 447836
rect 503126 447790 510866 447802
rect 503126 447378 510866 447390
rect 503126 447344 503138 447378
rect 510854 447344 510866 447378
rect 503126 447332 510866 447344
rect 503126 446920 510866 446932
rect 503126 446886 503138 446920
rect 510854 446886 510866 446920
rect 503126 446874 510866 446886
rect 503126 446462 510866 446474
rect 503126 446428 503138 446462
rect 510854 446428 510866 446462
rect 503126 446416 510866 446428
rect 503126 446004 510866 446016
rect 503126 445970 503138 446004
rect 510854 445970 510866 446004
rect 503126 445958 510866 445970
rect 503126 445546 510866 445558
rect 503126 445512 503138 445546
rect 510854 445512 510866 445546
rect 503126 445500 510866 445512
rect 503126 445088 510866 445100
rect 503126 445054 503138 445088
rect 510854 445054 510866 445088
rect 503126 445042 510866 445054
rect 503126 444630 510866 444642
rect 503126 444596 503138 444630
rect 510854 444596 510866 444630
rect 503126 444584 510866 444596
rect 503126 444172 510866 444184
rect 503126 444138 503138 444172
rect 510854 444138 510866 444172
rect 503126 444126 510866 444138
rect 503126 443714 510866 443726
rect 503126 443680 503138 443714
rect 510854 443680 510866 443714
rect 503126 443668 510866 443680
rect 503126 443256 510866 443268
rect 503126 443222 503138 443256
rect 510854 443222 510866 443256
rect 503126 443210 510866 443222
rect 503674 438124 504354 438178
rect 503674 438090 503728 438124
rect 503762 438090 503818 438124
rect 503852 438090 503908 438124
rect 503942 438090 503998 438124
rect 504032 438090 504088 438124
rect 504122 438090 504178 438124
rect 504212 438090 504268 438124
rect 504302 438090 504354 438124
rect 503674 438034 504354 438090
rect 503674 438000 503728 438034
rect 503762 438000 503818 438034
rect 503852 438000 503908 438034
rect 503942 438000 503998 438034
rect 504032 438000 504088 438034
rect 504122 438000 504178 438034
rect 504212 438000 504268 438034
rect 504302 438000 504354 438034
rect 503674 437944 504354 438000
rect 503674 437910 503728 437944
rect 503762 437910 503818 437944
rect 503852 437910 503908 437944
rect 503942 437910 503998 437944
rect 504032 437910 504088 437944
rect 504122 437910 504178 437944
rect 504212 437910 504268 437944
rect 504302 437910 504354 437944
rect 503674 437854 504354 437910
rect 503674 437820 503728 437854
rect 503762 437820 503818 437854
rect 503852 437820 503908 437854
rect 503942 437820 503998 437854
rect 504032 437820 504088 437854
rect 504122 437820 504178 437854
rect 504212 437820 504268 437854
rect 504302 437820 504354 437854
rect 503674 437764 504354 437820
rect 503674 437730 503728 437764
rect 503762 437730 503818 437764
rect 503852 437730 503908 437764
rect 503942 437730 503998 437764
rect 504032 437730 504088 437764
rect 504122 437730 504178 437764
rect 504212 437730 504268 437764
rect 504302 437730 504354 437764
rect 503674 437674 504354 437730
rect 503674 437640 503728 437674
rect 503762 437640 503818 437674
rect 503852 437640 503908 437674
rect 503942 437640 503998 437674
rect 504032 437640 504088 437674
rect 504122 437640 504178 437674
rect 504212 437640 504268 437674
rect 504302 437640 504354 437674
rect 503674 437584 504354 437640
rect 503674 437550 503728 437584
rect 503762 437550 503818 437584
rect 503852 437550 503908 437584
rect 503942 437550 503998 437584
rect 504032 437550 504088 437584
rect 504122 437550 504178 437584
rect 504212 437550 504268 437584
rect 504302 437550 504354 437584
rect 503674 437498 504354 437550
rect 504962 438124 505642 438178
rect 504962 438090 505016 438124
rect 505050 438090 505106 438124
rect 505140 438090 505196 438124
rect 505230 438090 505286 438124
rect 505320 438090 505376 438124
rect 505410 438090 505466 438124
rect 505500 438090 505556 438124
rect 505590 438090 505642 438124
rect 504962 438034 505642 438090
rect 504962 438000 505016 438034
rect 505050 438000 505106 438034
rect 505140 438000 505196 438034
rect 505230 438000 505286 438034
rect 505320 438000 505376 438034
rect 505410 438000 505466 438034
rect 505500 438000 505556 438034
rect 505590 438000 505642 438034
rect 504962 437944 505642 438000
rect 504962 437910 505016 437944
rect 505050 437910 505106 437944
rect 505140 437910 505196 437944
rect 505230 437910 505286 437944
rect 505320 437910 505376 437944
rect 505410 437910 505466 437944
rect 505500 437910 505556 437944
rect 505590 437910 505642 437944
rect 504962 437854 505642 437910
rect 504962 437820 505016 437854
rect 505050 437820 505106 437854
rect 505140 437820 505196 437854
rect 505230 437820 505286 437854
rect 505320 437820 505376 437854
rect 505410 437820 505466 437854
rect 505500 437820 505556 437854
rect 505590 437820 505642 437854
rect 504962 437764 505642 437820
rect 504962 437730 505016 437764
rect 505050 437730 505106 437764
rect 505140 437730 505196 437764
rect 505230 437730 505286 437764
rect 505320 437730 505376 437764
rect 505410 437730 505466 437764
rect 505500 437730 505556 437764
rect 505590 437730 505642 437764
rect 504962 437674 505642 437730
rect 504962 437640 505016 437674
rect 505050 437640 505106 437674
rect 505140 437640 505196 437674
rect 505230 437640 505286 437674
rect 505320 437640 505376 437674
rect 505410 437640 505466 437674
rect 505500 437640 505556 437674
rect 505590 437640 505642 437674
rect 504962 437584 505642 437640
rect 504962 437550 505016 437584
rect 505050 437550 505106 437584
rect 505140 437550 505196 437584
rect 505230 437550 505286 437584
rect 505320 437550 505376 437584
rect 505410 437550 505466 437584
rect 505500 437550 505556 437584
rect 505590 437550 505642 437584
rect 504962 437498 505642 437550
rect 506250 438124 506930 438178
rect 506250 438090 506304 438124
rect 506338 438090 506394 438124
rect 506428 438090 506484 438124
rect 506518 438090 506574 438124
rect 506608 438090 506664 438124
rect 506698 438090 506754 438124
rect 506788 438090 506844 438124
rect 506878 438090 506930 438124
rect 506250 438034 506930 438090
rect 506250 438000 506304 438034
rect 506338 438000 506394 438034
rect 506428 438000 506484 438034
rect 506518 438000 506574 438034
rect 506608 438000 506664 438034
rect 506698 438000 506754 438034
rect 506788 438000 506844 438034
rect 506878 438000 506930 438034
rect 506250 437944 506930 438000
rect 506250 437910 506304 437944
rect 506338 437910 506394 437944
rect 506428 437910 506484 437944
rect 506518 437910 506574 437944
rect 506608 437910 506664 437944
rect 506698 437910 506754 437944
rect 506788 437910 506844 437944
rect 506878 437910 506930 437944
rect 506250 437854 506930 437910
rect 506250 437820 506304 437854
rect 506338 437820 506394 437854
rect 506428 437820 506484 437854
rect 506518 437820 506574 437854
rect 506608 437820 506664 437854
rect 506698 437820 506754 437854
rect 506788 437820 506844 437854
rect 506878 437820 506930 437854
rect 506250 437764 506930 437820
rect 506250 437730 506304 437764
rect 506338 437730 506394 437764
rect 506428 437730 506484 437764
rect 506518 437730 506574 437764
rect 506608 437730 506664 437764
rect 506698 437730 506754 437764
rect 506788 437730 506844 437764
rect 506878 437730 506930 437764
rect 506250 437674 506930 437730
rect 506250 437640 506304 437674
rect 506338 437640 506394 437674
rect 506428 437640 506484 437674
rect 506518 437640 506574 437674
rect 506608 437640 506664 437674
rect 506698 437640 506754 437674
rect 506788 437640 506844 437674
rect 506878 437640 506930 437674
rect 506250 437584 506930 437640
rect 506250 437550 506304 437584
rect 506338 437550 506394 437584
rect 506428 437550 506484 437584
rect 506518 437550 506574 437584
rect 506608 437550 506664 437584
rect 506698 437550 506754 437584
rect 506788 437550 506844 437584
rect 506878 437550 506930 437584
rect 506250 437498 506930 437550
rect 507538 438124 508218 438178
rect 507538 438090 507592 438124
rect 507626 438090 507682 438124
rect 507716 438090 507772 438124
rect 507806 438090 507862 438124
rect 507896 438090 507952 438124
rect 507986 438090 508042 438124
rect 508076 438090 508132 438124
rect 508166 438090 508218 438124
rect 507538 438034 508218 438090
rect 507538 438000 507592 438034
rect 507626 438000 507682 438034
rect 507716 438000 507772 438034
rect 507806 438000 507862 438034
rect 507896 438000 507952 438034
rect 507986 438000 508042 438034
rect 508076 438000 508132 438034
rect 508166 438000 508218 438034
rect 507538 437944 508218 438000
rect 507538 437910 507592 437944
rect 507626 437910 507682 437944
rect 507716 437910 507772 437944
rect 507806 437910 507862 437944
rect 507896 437910 507952 437944
rect 507986 437910 508042 437944
rect 508076 437910 508132 437944
rect 508166 437910 508218 437944
rect 507538 437854 508218 437910
rect 507538 437820 507592 437854
rect 507626 437820 507682 437854
rect 507716 437820 507772 437854
rect 507806 437820 507862 437854
rect 507896 437820 507952 437854
rect 507986 437820 508042 437854
rect 508076 437820 508132 437854
rect 508166 437820 508218 437854
rect 507538 437764 508218 437820
rect 507538 437730 507592 437764
rect 507626 437730 507682 437764
rect 507716 437730 507772 437764
rect 507806 437730 507862 437764
rect 507896 437730 507952 437764
rect 507986 437730 508042 437764
rect 508076 437730 508132 437764
rect 508166 437730 508218 437764
rect 507538 437674 508218 437730
rect 507538 437640 507592 437674
rect 507626 437640 507682 437674
rect 507716 437640 507772 437674
rect 507806 437640 507862 437674
rect 507896 437640 507952 437674
rect 507986 437640 508042 437674
rect 508076 437640 508132 437674
rect 508166 437640 508218 437674
rect 507538 437584 508218 437640
rect 507538 437550 507592 437584
rect 507626 437550 507682 437584
rect 507716 437550 507772 437584
rect 507806 437550 507862 437584
rect 507896 437550 507952 437584
rect 507986 437550 508042 437584
rect 508076 437550 508132 437584
rect 508166 437550 508218 437584
rect 507538 437498 508218 437550
rect 508826 438124 509506 438178
rect 508826 438090 508880 438124
rect 508914 438090 508970 438124
rect 509004 438090 509060 438124
rect 509094 438090 509150 438124
rect 509184 438090 509240 438124
rect 509274 438090 509330 438124
rect 509364 438090 509420 438124
rect 509454 438090 509506 438124
rect 508826 438034 509506 438090
rect 508826 438000 508880 438034
rect 508914 438000 508970 438034
rect 509004 438000 509060 438034
rect 509094 438000 509150 438034
rect 509184 438000 509240 438034
rect 509274 438000 509330 438034
rect 509364 438000 509420 438034
rect 509454 438000 509506 438034
rect 508826 437944 509506 438000
rect 508826 437910 508880 437944
rect 508914 437910 508970 437944
rect 509004 437910 509060 437944
rect 509094 437910 509150 437944
rect 509184 437910 509240 437944
rect 509274 437910 509330 437944
rect 509364 437910 509420 437944
rect 509454 437910 509506 437944
rect 508826 437854 509506 437910
rect 508826 437820 508880 437854
rect 508914 437820 508970 437854
rect 509004 437820 509060 437854
rect 509094 437820 509150 437854
rect 509184 437820 509240 437854
rect 509274 437820 509330 437854
rect 509364 437820 509420 437854
rect 509454 437820 509506 437854
rect 508826 437764 509506 437820
rect 508826 437730 508880 437764
rect 508914 437730 508970 437764
rect 509004 437730 509060 437764
rect 509094 437730 509150 437764
rect 509184 437730 509240 437764
rect 509274 437730 509330 437764
rect 509364 437730 509420 437764
rect 509454 437730 509506 437764
rect 508826 437674 509506 437730
rect 508826 437640 508880 437674
rect 508914 437640 508970 437674
rect 509004 437640 509060 437674
rect 509094 437640 509150 437674
rect 509184 437640 509240 437674
rect 509274 437640 509330 437674
rect 509364 437640 509420 437674
rect 509454 437640 509506 437674
rect 508826 437584 509506 437640
rect 508826 437550 508880 437584
rect 508914 437550 508970 437584
rect 509004 437550 509060 437584
rect 509094 437550 509150 437584
rect 509184 437550 509240 437584
rect 509274 437550 509330 437584
rect 509364 437550 509420 437584
rect 509454 437550 509506 437584
rect 508826 437498 509506 437550
rect 510114 438124 510794 438178
rect 510114 438090 510168 438124
rect 510202 438090 510258 438124
rect 510292 438090 510348 438124
rect 510382 438090 510438 438124
rect 510472 438090 510528 438124
rect 510562 438090 510618 438124
rect 510652 438090 510708 438124
rect 510742 438090 510794 438124
rect 510114 438034 510794 438090
rect 510114 438000 510168 438034
rect 510202 438000 510258 438034
rect 510292 438000 510348 438034
rect 510382 438000 510438 438034
rect 510472 438000 510528 438034
rect 510562 438000 510618 438034
rect 510652 438000 510708 438034
rect 510742 438000 510794 438034
rect 510114 437944 510794 438000
rect 510114 437910 510168 437944
rect 510202 437910 510258 437944
rect 510292 437910 510348 437944
rect 510382 437910 510438 437944
rect 510472 437910 510528 437944
rect 510562 437910 510618 437944
rect 510652 437910 510708 437944
rect 510742 437910 510794 437944
rect 510114 437854 510794 437910
rect 510114 437820 510168 437854
rect 510202 437820 510258 437854
rect 510292 437820 510348 437854
rect 510382 437820 510438 437854
rect 510472 437820 510528 437854
rect 510562 437820 510618 437854
rect 510652 437820 510708 437854
rect 510742 437820 510794 437854
rect 510114 437764 510794 437820
rect 510114 437730 510168 437764
rect 510202 437730 510258 437764
rect 510292 437730 510348 437764
rect 510382 437730 510438 437764
rect 510472 437730 510528 437764
rect 510562 437730 510618 437764
rect 510652 437730 510708 437764
rect 510742 437730 510794 437764
rect 510114 437674 510794 437730
rect 510114 437640 510168 437674
rect 510202 437640 510258 437674
rect 510292 437640 510348 437674
rect 510382 437640 510438 437674
rect 510472 437640 510528 437674
rect 510562 437640 510618 437674
rect 510652 437640 510708 437674
rect 510742 437640 510794 437674
rect 510114 437584 510794 437640
rect 510114 437550 510168 437584
rect 510202 437550 510258 437584
rect 510292 437550 510348 437584
rect 510382 437550 510438 437584
rect 510472 437550 510528 437584
rect 510562 437550 510618 437584
rect 510652 437550 510708 437584
rect 510742 437550 510794 437584
rect 510114 437498 510794 437550
rect 511402 438124 512082 438178
rect 511402 438090 511456 438124
rect 511490 438090 511546 438124
rect 511580 438090 511636 438124
rect 511670 438090 511726 438124
rect 511760 438090 511816 438124
rect 511850 438090 511906 438124
rect 511940 438090 511996 438124
rect 512030 438090 512082 438124
rect 511402 438034 512082 438090
rect 511402 438000 511456 438034
rect 511490 438000 511546 438034
rect 511580 438000 511636 438034
rect 511670 438000 511726 438034
rect 511760 438000 511816 438034
rect 511850 438000 511906 438034
rect 511940 438000 511996 438034
rect 512030 438000 512082 438034
rect 511402 437944 512082 438000
rect 511402 437910 511456 437944
rect 511490 437910 511546 437944
rect 511580 437910 511636 437944
rect 511670 437910 511726 437944
rect 511760 437910 511816 437944
rect 511850 437910 511906 437944
rect 511940 437910 511996 437944
rect 512030 437910 512082 437944
rect 511402 437854 512082 437910
rect 511402 437820 511456 437854
rect 511490 437820 511546 437854
rect 511580 437820 511636 437854
rect 511670 437820 511726 437854
rect 511760 437820 511816 437854
rect 511850 437820 511906 437854
rect 511940 437820 511996 437854
rect 512030 437820 512082 437854
rect 511402 437764 512082 437820
rect 511402 437730 511456 437764
rect 511490 437730 511546 437764
rect 511580 437730 511636 437764
rect 511670 437730 511726 437764
rect 511760 437730 511816 437764
rect 511850 437730 511906 437764
rect 511940 437730 511996 437764
rect 512030 437730 512082 437764
rect 511402 437674 512082 437730
rect 511402 437640 511456 437674
rect 511490 437640 511546 437674
rect 511580 437640 511636 437674
rect 511670 437640 511726 437674
rect 511760 437640 511816 437674
rect 511850 437640 511906 437674
rect 511940 437640 511996 437674
rect 512030 437640 512082 437674
rect 511402 437584 512082 437640
rect 511402 437550 511456 437584
rect 511490 437550 511546 437584
rect 511580 437550 511636 437584
rect 511670 437550 511726 437584
rect 511760 437550 511816 437584
rect 511850 437550 511906 437584
rect 511940 437550 511996 437584
rect 512030 437550 512082 437584
rect 511402 437498 512082 437550
rect 512690 438124 513370 438178
rect 512690 438090 512744 438124
rect 512778 438090 512834 438124
rect 512868 438090 512924 438124
rect 512958 438090 513014 438124
rect 513048 438090 513104 438124
rect 513138 438090 513194 438124
rect 513228 438090 513284 438124
rect 513318 438090 513370 438124
rect 512690 438034 513370 438090
rect 512690 438000 512744 438034
rect 512778 438000 512834 438034
rect 512868 438000 512924 438034
rect 512958 438000 513014 438034
rect 513048 438000 513104 438034
rect 513138 438000 513194 438034
rect 513228 438000 513284 438034
rect 513318 438000 513370 438034
rect 512690 437944 513370 438000
rect 512690 437910 512744 437944
rect 512778 437910 512834 437944
rect 512868 437910 512924 437944
rect 512958 437910 513014 437944
rect 513048 437910 513104 437944
rect 513138 437910 513194 437944
rect 513228 437910 513284 437944
rect 513318 437910 513370 437944
rect 512690 437854 513370 437910
rect 512690 437820 512744 437854
rect 512778 437820 512834 437854
rect 512868 437820 512924 437854
rect 512958 437820 513014 437854
rect 513048 437820 513104 437854
rect 513138 437820 513194 437854
rect 513228 437820 513284 437854
rect 513318 437820 513370 437854
rect 512690 437764 513370 437820
rect 512690 437730 512744 437764
rect 512778 437730 512834 437764
rect 512868 437730 512924 437764
rect 512958 437730 513014 437764
rect 513048 437730 513104 437764
rect 513138 437730 513194 437764
rect 513228 437730 513284 437764
rect 513318 437730 513370 437764
rect 512690 437674 513370 437730
rect 512690 437640 512744 437674
rect 512778 437640 512834 437674
rect 512868 437640 512924 437674
rect 512958 437640 513014 437674
rect 513048 437640 513104 437674
rect 513138 437640 513194 437674
rect 513228 437640 513284 437674
rect 513318 437640 513370 437674
rect 512690 437584 513370 437640
rect 512690 437550 512744 437584
rect 512778 437550 512834 437584
rect 512868 437550 512924 437584
rect 512958 437550 513014 437584
rect 513048 437550 513104 437584
rect 513138 437550 513194 437584
rect 513228 437550 513284 437584
rect 513318 437550 513370 437584
rect 512690 437498 513370 437550
rect 503674 436836 504354 436890
rect 503674 436802 503728 436836
rect 503762 436802 503818 436836
rect 503852 436802 503908 436836
rect 503942 436802 503998 436836
rect 504032 436802 504088 436836
rect 504122 436802 504178 436836
rect 504212 436802 504268 436836
rect 504302 436802 504354 436836
rect 503674 436746 504354 436802
rect 503674 436712 503728 436746
rect 503762 436712 503818 436746
rect 503852 436712 503908 436746
rect 503942 436712 503998 436746
rect 504032 436712 504088 436746
rect 504122 436712 504178 436746
rect 504212 436712 504268 436746
rect 504302 436712 504354 436746
rect 503674 436656 504354 436712
rect 503674 436622 503728 436656
rect 503762 436622 503818 436656
rect 503852 436622 503908 436656
rect 503942 436622 503998 436656
rect 504032 436622 504088 436656
rect 504122 436622 504178 436656
rect 504212 436622 504268 436656
rect 504302 436622 504354 436656
rect 503674 436566 504354 436622
rect 503674 436532 503728 436566
rect 503762 436532 503818 436566
rect 503852 436532 503908 436566
rect 503942 436532 503998 436566
rect 504032 436532 504088 436566
rect 504122 436532 504178 436566
rect 504212 436532 504268 436566
rect 504302 436532 504354 436566
rect 503674 436476 504354 436532
rect 503674 436442 503728 436476
rect 503762 436442 503818 436476
rect 503852 436442 503908 436476
rect 503942 436442 503998 436476
rect 504032 436442 504088 436476
rect 504122 436442 504178 436476
rect 504212 436442 504268 436476
rect 504302 436442 504354 436476
rect 503674 436386 504354 436442
rect 503674 436352 503728 436386
rect 503762 436352 503818 436386
rect 503852 436352 503908 436386
rect 503942 436352 503998 436386
rect 504032 436352 504088 436386
rect 504122 436352 504178 436386
rect 504212 436352 504268 436386
rect 504302 436352 504354 436386
rect 503674 436296 504354 436352
rect 503674 436262 503728 436296
rect 503762 436262 503818 436296
rect 503852 436262 503908 436296
rect 503942 436262 503998 436296
rect 504032 436262 504088 436296
rect 504122 436262 504178 436296
rect 504212 436262 504268 436296
rect 504302 436262 504354 436296
rect 503674 436210 504354 436262
rect 504962 436836 505642 436890
rect 504962 436802 505016 436836
rect 505050 436802 505106 436836
rect 505140 436802 505196 436836
rect 505230 436802 505286 436836
rect 505320 436802 505376 436836
rect 505410 436802 505466 436836
rect 505500 436802 505556 436836
rect 505590 436802 505642 436836
rect 504962 436746 505642 436802
rect 504962 436712 505016 436746
rect 505050 436712 505106 436746
rect 505140 436712 505196 436746
rect 505230 436712 505286 436746
rect 505320 436712 505376 436746
rect 505410 436712 505466 436746
rect 505500 436712 505556 436746
rect 505590 436712 505642 436746
rect 504962 436656 505642 436712
rect 504962 436622 505016 436656
rect 505050 436622 505106 436656
rect 505140 436622 505196 436656
rect 505230 436622 505286 436656
rect 505320 436622 505376 436656
rect 505410 436622 505466 436656
rect 505500 436622 505556 436656
rect 505590 436622 505642 436656
rect 504962 436566 505642 436622
rect 504962 436532 505016 436566
rect 505050 436532 505106 436566
rect 505140 436532 505196 436566
rect 505230 436532 505286 436566
rect 505320 436532 505376 436566
rect 505410 436532 505466 436566
rect 505500 436532 505556 436566
rect 505590 436532 505642 436566
rect 504962 436476 505642 436532
rect 504962 436442 505016 436476
rect 505050 436442 505106 436476
rect 505140 436442 505196 436476
rect 505230 436442 505286 436476
rect 505320 436442 505376 436476
rect 505410 436442 505466 436476
rect 505500 436442 505556 436476
rect 505590 436442 505642 436476
rect 504962 436386 505642 436442
rect 504962 436352 505016 436386
rect 505050 436352 505106 436386
rect 505140 436352 505196 436386
rect 505230 436352 505286 436386
rect 505320 436352 505376 436386
rect 505410 436352 505466 436386
rect 505500 436352 505556 436386
rect 505590 436352 505642 436386
rect 504962 436296 505642 436352
rect 504962 436262 505016 436296
rect 505050 436262 505106 436296
rect 505140 436262 505196 436296
rect 505230 436262 505286 436296
rect 505320 436262 505376 436296
rect 505410 436262 505466 436296
rect 505500 436262 505556 436296
rect 505590 436262 505642 436296
rect 504962 436210 505642 436262
rect 506250 436836 506930 436890
rect 506250 436802 506304 436836
rect 506338 436802 506394 436836
rect 506428 436802 506484 436836
rect 506518 436802 506574 436836
rect 506608 436802 506664 436836
rect 506698 436802 506754 436836
rect 506788 436802 506844 436836
rect 506878 436802 506930 436836
rect 506250 436746 506930 436802
rect 506250 436712 506304 436746
rect 506338 436712 506394 436746
rect 506428 436712 506484 436746
rect 506518 436712 506574 436746
rect 506608 436712 506664 436746
rect 506698 436712 506754 436746
rect 506788 436712 506844 436746
rect 506878 436712 506930 436746
rect 506250 436656 506930 436712
rect 506250 436622 506304 436656
rect 506338 436622 506394 436656
rect 506428 436622 506484 436656
rect 506518 436622 506574 436656
rect 506608 436622 506664 436656
rect 506698 436622 506754 436656
rect 506788 436622 506844 436656
rect 506878 436622 506930 436656
rect 506250 436566 506930 436622
rect 506250 436532 506304 436566
rect 506338 436532 506394 436566
rect 506428 436532 506484 436566
rect 506518 436532 506574 436566
rect 506608 436532 506664 436566
rect 506698 436532 506754 436566
rect 506788 436532 506844 436566
rect 506878 436532 506930 436566
rect 506250 436476 506930 436532
rect 506250 436442 506304 436476
rect 506338 436442 506394 436476
rect 506428 436442 506484 436476
rect 506518 436442 506574 436476
rect 506608 436442 506664 436476
rect 506698 436442 506754 436476
rect 506788 436442 506844 436476
rect 506878 436442 506930 436476
rect 506250 436386 506930 436442
rect 506250 436352 506304 436386
rect 506338 436352 506394 436386
rect 506428 436352 506484 436386
rect 506518 436352 506574 436386
rect 506608 436352 506664 436386
rect 506698 436352 506754 436386
rect 506788 436352 506844 436386
rect 506878 436352 506930 436386
rect 506250 436296 506930 436352
rect 506250 436262 506304 436296
rect 506338 436262 506394 436296
rect 506428 436262 506484 436296
rect 506518 436262 506574 436296
rect 506608 436262 506664 436296
rect 506698 436262 506754 436296
rect 506788 436262 506844 436296
rect 506878 436262 506930 436296
rect 506250 436210 506930 436262
rect 507538 436836 508218 436890
rect 507538 436802 507592 436836
rect 507626 436802 507682 436836
rect 507716 436802 507772 436836
rect 507806 436802 507862 436836
rect 507896 436802 507952 436836
rect 507986 436802 508042 436836
rect 508076 436802 508132 436836
rect 508166 436802 508218 436836
rect 507538 436746 508218 436802
rect 507538 436712 507592 436746
rect 507626 436712 507682 436746
rect 507716 436712 507772 436746
rect 507806 436712 507862 436746
rect 507896 436712 507952 436746
rect 507986 436712 508042 436746
rect 508076 436712 508132 436746
rect 508166 436712 508218 436746
rect 507538 436656 508218 436712
rect 507538 436622 507592 436656
rect 507626 436622 507682 436656
rect 507716 436622 507772 436656
rect 507806 436622 507862 436656
rect 507896 436622 507952 436656
rect 507986 436622 508042 436656
rect 508076 436622 508132 436656
rect 508166 436622 508218 436656
rect 507538 436566 508218 436622
rect 507538 436532 507592 436566
rect 507626 436532 507682 436566
rect 507716 436532 507772 436566
rect 507806 436532 507862 436566
rect 507896 436532 507952 436566
rect 507986 436532 508042 436566
rect 508076 436532 508132 436566
rect 508166 436532 508218 436566
rect 507538 436476 508218 436532
rect 507538 436442 507592 436476
rect 507626 436442 507682 436476
rect 507716 436442 507772 436476
rect 507806 436442 507862 436476
rect 507896 436442 507952 436476
rect 507986 436442 508042 436476
rect 508076 436442 508132 436476
rect 508166 436442 508218 436476
rect 507538 436386 508218 436442
rect 507538 436352 507592 436386
rect 507626 436352 507682 436386
rect 507716 436352 507772 436386
rect 507806 436352 507862 436386
rect 507896 436352 507952 436386
rect 507986 436352 508042 436386
rect 508076 436352 508132 436386
rect 508166 436352 508218 436386
rect 507538 436296 508218 436352
rect 507538 436262 507592 436296
rect 507626 436262 507682 436296
rect 507716 436262 507772 436296
rect 507806 436262 507862 436296
rect 507896 436262 507952 436296
rect 507986 436262 508042 436296
rect 508076 436262 508132 436296
rect 508166 436262 508218 436296
rect 507538 436210 508218 436262
rect 508826 436836 509506 436890
rect 508826 436802 508880 436836
rect 508914 436802 508970 436836
rect 509004 436802 509060 436836
rect 509094 436802 509150 436836
rect 509184 436802 509240 436836
rect 509274 436802 509330 436836
rect 509364 436802 509420 436836
rect 509454 436802 509506 436836
rect 508826 436746 509506 436802
rect 508826 436712 508880 436746
rect 508914 436712 508970 436746
rect 509004 436712 509060 436746
rect 509094 436712 509150 436746
rect 509184 436712 509240 436746
rect 509274 436712 509330 436746
rect 509364 436712 509420 436746
rect 509454 436712 509506 436746
rect 508826 436656 509506 436712
rect 508826 436622 508880 436656
rect 508914 436622 508970 436656
rect 509004 436622 509060 436656
rect 509094 436622 509150 436656
rect 509184 436622 509240 436656
rect 509274 436622 509330 436656
rect 509364 436622 509420 436656
rect 509454 436622 509506 436656
rect 508826 436566 509506 436622
rect 508826 436532 508880 436566
rect 508914 436532 508970 436566
rect 509004 436532 509060 436566
rect 509094 436532 509150 436566
rect 509184 436532 509240 436566
rect 509274 436532 509330 436566
rect 509364 436532 509420 436566
rect 509454 436532 509506 436566
rect 508826 436476 509506 436532
rect 508826 436442 508880 436476
rect 508914 436442 508970 436476
rect 509004 436442 509060 436476
rect 509094 436442 509150 436476
rect 509184 436442 509240 436476
rect 509274 436442 509330 436476
rect 509364 436442 509420 436476
rect 509454 436442 509506 436476
rect 508826 436386 509506 436442
rect 508826 436352 508880 436386
rect 508914 436352 508970 436386
rect 509004 436352 509060 436386
rect 509094 436352 509150 436386
rect 509184 436352 509240 436386
rect 509274 436352 509330 436386
rect 509364 436352 509420 436386
rect 509454 436352 509506 436386
rect 508826 436296 509506 436352
rect 508826 436262 508880 436296
rect 508914 436262 508970 436296
rect 509004 436262 509060 436296
rect 509094 436262 509150 436296
rect 509184 436262 509240 436296
rect 509274 436262 509330 436296
rect 509364 436262 509420 436296
rect 509454 436262 509506 436296
rect 508826 436210 509506 436262
rect 510114 436836 510794 436890
rect 510114 436802 510168 436836
rect 510202 436802 510258 436836
rect 510292 436802 510348 436836
rect 510382 436802 510438 436836
rect 510472 436802 510528 436836
rect 510562 436802 510618 436836
rect 510652 436802 510708 436836
rect 510742 436802 510794 436836
rect 510114 436746 510794 436802
rect 510114 436712 510168 436746
rect 510202 436712 510258 436746
rect 510292 436712 510348 436746
rect 510382 436712 510438 436746
rect 510472 436712 510528 436746
rect 510562 436712 510618 436746
rect 510652 436712 510708 436746
rect 510742 436712 510794 436746
rect 510114 436656 510794 436712
rect 510114 436622 510168 436656
rect 510202 436622 510258 436656
rect 510292 436622 510348 436656
rect 510382 436622 510438 436656
rect 510472 436622 510528 436656
rect 510562 436622 510618 436656
rect 510652 436622 510708 436656
rect 510742 436622 510794 436656
rect 510114 436566 510794 436622
rect 510114 436532 510168 436566
rect 510202 436532 510258 436566
rect 510292 436532 510348 436566
rect 510382 436532 510438 436566
rect 510472 436532 510528 436566
rect 510562 436532 510618 436566
rect 510652 436532 510708 436566
rect 510742 436532 510794 436566
rect 510114 436476 510794 436532
rect 510114 436442 510168 436476
rect 510202 436442 510258 436476
rect 510292 436442 510348 436476
rect 510382 436442 510438 436476
rect 510472 436442 510528 436476
rect 510562 436442 510618 436476
rect 510652 436442 510708 436476
rect 510742 436442 510794 436476
rect 510114 436386 510794 436442
rect 510114 436352 510168 436386
rect 510202 436352 510258 436386
rect 510292 436352 510348 436386
rect 510382 436352 510438 436386
rect 510472 436352 510528 436386
rect 510562 436352 510618 436386
rect 510652 436352 510708 436386
rect 510742 436352 510794 436386
rect 510114 436296 510794 436352
rect 510114 436262 510168 436296
rect 510202 436262 510258 436296
rect 510292 436262 510348 436296
rect 510382 436262 510438 436296
rect 510472 436262 510528 436296
rect 510562 436262 510618 436296
rect 510652 436262 510708 436296
rect 510742 436262 510794 436296
rect 510114 436210 510794 436262
rect 511402 436836 512082 436890
rect 511402 436802 511456 436836
rect 511490 436802 511546 436836
rect 511580 436802 511636 436836
rect 511670 436802 511726 436836
rect 511760 436802 511816 436836
rect 511850 436802 511906 436836
rect 511940 436802 511996 436836
rect 512030 436802 512082 436836
rect 511402 436746 512082 436802
rect 511402 436712 511456 436746
rect 511490 436712 511546 436746
rect 511580 436712 511636 436746
rect 511670 436712 511726 436746
rect 511760 436712 511816 436746
rect 511850 436712 511906 436746
rect 511940 436712 511996 436746
rect 512030 436712 512082 436746
rect 511402 436656 512082 436712
rect 511402 436622 511456 436656
rect 511490 436622 511546 436656
rect 511580 436622 511636 436656
rect 511670 436622 511726 436656
rect 511760 436622 511816 436656
rect 511850 436622 511906 436656
rect 511940 436622 511996 436656
rect 512030 436622 512082 436656
rect 511402 436566 512082 436622
rect 511402 436532 511456 436566
rect 511490 436532 511546 436566
rect 511580 436532 511636 436566
rect 511670 436532 511726 436566
rect 511760 436532 511816 436566
rect 511850 436532 511906 436566
rect 511940 436532 511996 436566
rect 512030 436532 512082 436566
rect 511402 436476 512082 436532
rect 511402 436442 511456 436476
rect 511490 436442 511546 436476
rect 511580 436442 511636 436476
rect 511670 436442 511726 436476
rect 511760 436442 511816 436476
rect 511850 436442 511906 436476
rect 511940 436442 511996 436476
rect 512030 436442 512082 436476
rect 511402 436386 512082 436442
rect 511402 436352 511456 436386
rect 511490 436352 511546 436386
rect 511580 436352 511636 436386
rect 511670 436352 511726 436386
rect 511760 436352 511816 436386
rect 511850 436352 511906 436386
rect 511940 436352 511996 436386
rect 512030 436352 512082 436386
rect 511402 436296 512082 436352
rect 511402 436262 511456 436296
rect 511490 436262 511546 436296
rect 511580 436262 511636 436296
rect 511670 436262 511726 436296
rect 511760 436262 511816 436296
rect 511850 436262 511906 436296
rect 511940 436262 511996 436296
rect 512030 436262 512082 436296
rect 511402 436210 512082 436262
rect 512690 436836 513370 436890
rect 512690 436802 512744 436836
rect 512778 436802 512834 436836
rect 512868 436802 512924 436836
rect 512958 436802 513014 436836
rect 513048 436802 513104 436836
rect 513138 436802 513194 436836
rect 513228 436802 513284 436836
rect 513318 436802 513370 436836
rect 512690 436746 513370 436802
rect 512690 436712 512744 436746
rect 512778 436712 512834 436746
rect 512868 436712 512924 436746
rect 512958 436712 513014 436746
rect 513048 436712 513104 436746
rect 513138 436712 513194 436746
rect 513228 436712 513284 436746
rect 513318 436712 513370 436746
rect 512690 436656 513370 436712
rect 512690 436622 512744 436656
rect 512778 436622 512834 436656
rect 512868 436622 512924 436656
rect 512958 436622 513014 436656
rect 513048 436622 513104 436656
rect 513138 436622 513194 436656
rect 513228 436622 513284 436656
rect 513318 436622 513370 436656
rect 512690 436566 513370 436622
rect 512690 436532 512744 436566
rect 512778 436532 512834 436566
rect 512868 436532 512924 436566
rect 512958 436532 513014 436566
rect 513048 436532 513104 436566
rect 513138 436532 513194 436566
rect 513228 436532 513284 436566
rect 513318 436532 513370 436566
rect 512690 436476 513370 436532
rect 512690 436442 512744 436476
rect 512778 436442 512834 436476
rect 512868 436442 512924 436476
rect 512958 436442 513014 436476
rect 513048 436442 513104 436476
rect 513138 436442 513194 436476
rect 513228 436442 513284 436476
rect 513318 436442 513370 436476
rect 512690 436386 513370 436442
rect 512690 436352 512744 436386
rect 512778 436352 512834 436386
rect 512868 436352 512924 436386
rect 512958 436352 513014 436386
rect 513048 436352 513104 436386
rect 513138 436352 513194 436386
rect 513228 436352 513284 436386
rect 513318 436352 513370 436386
rect 512690 436296 513370 436352
rect 512690 436262 512744 436296
rect 512778 436262 512834 436296
rect 512868 436262 512924 436296
rect 512958 436262 513014 436296
rect 513048 436262 513104 436296
rect 513138 436262 513194 436296
rect 513228 436262 513284 436296
rect 513318 436262 513370 436296
rect 512690 436210 513370 436262
rect 503674 435548 504354 435602
rect 503674 435514 503728 435548
rect 503762 435514 503818 435548
rect 503852 435514 503908 435548
rect 503942 435514 503998 435548
rect 504032 435514 504088 435548
rect 504122 435514 504178 435548
rect 504212 435514 504268 435548
rect 504302 435514 504354 435548
rect 503674 435458 504354 435514
rect 503674 435424 503728 435458
rect 503762 435424 503818 435458
rect 503852 435424 503908 435458
rect 503942 435424 503998 435458
rect 504032 435424 504088 435458
rect 504122 435424 504178 435458
rect 504212 435424 504268 435458
rect 504302 435424 504354 435458
rect 503674 435368 504354 435424
rect 503674 435334 503728 435368
rect 503762 435334 503818 435368
rect 503852 435334 503908 435368
rect 503942 435334 503998 435368
rect 504032 435334 504088 435368
rect 504122 435334 504178 435368
rect 504212 435334 504268 435368
rect 504302 435334 504354 435368
rect 503674 435278 504354 435334
rect 503674 435244 503728 435278
rect 503762 435244 503818 435278
rect 503852 435244 503908 435278
rect 503942 435244 503998 435278
rect 504032 435244 504088 435278
rect 504122 435244 504178 435278
rect 504212 435244 504268 435278
rect 504302 435244 504354 435278
rect 503674 435188 504354 435244
rect 503674 435154 503728 435188
rect 503762 435154 503818 435188
rect 503852 435154 503908 435188
rect 503942 435154 503998 435188
rect 504032 435154 504088 435188
rect 504122 435154 504178 435188
rect 504212 435154 504268 435188
rect 504302 435154 504354 435188
rect 503674 435098 504354 435154
rect 503674 435064 503728 435098
rect 503762 435064 503818 435098
rect 503852 435064 503908 435098
rect 503942 435064 503998 435098
rect 504032 435064 504088 435098
rect 504122 435064 504178 435098
rect 504212 435064 504268 435098
rect 504302 435064 504354 435098
rect 503674 435008 504354 435064
rect 503674 434974 503728 435008
rect 503762 434974 503818 435008
rect 503852 434974 503908 435008
rect 503942 434974 503998 435008
rect 504032 434974 504088 435008
rect 504122 434974 504178 435008
rect 504212 434974 504268 435008
rect 504302 434974 504354 435008
rect 503674 434922 504354 434974
rect 504962 435548 505642 435602
rect 504962 435514 505016 435548
rect 505050 435514 505106 435548
rect 505140 435514 505196 435548
rect 505230 435514 505286 435548
rect 505320 435514 505376 435548
rect 505410 435514 505466 435548
rect 505500 435514 505556 435548
rect 505590 435514 505642 435548
rect 504962 435458 505642 435514
rect 504962 435424 505016 435458
rect 505050 435424 505106 435458
rect 505140 435424 505196 435458
rect 505230 435424 505286 435458
rect 505320 435424 505376 435458
rect 505410 435424 505466 435458
rect 505500 435424 505556 435458
rect 505590 435424 505642 435458
rect 504962 435368 505642 435424
rect 504962 435334 505016 435368
rect 505050 435334 505106 435368
rect 505140 435334 505196 435368
rect 505230 435334 505286 435368
rect 505320 435334 505376 435368
rect 505410 435334 505466 435368
rect 505500 435334 505556 435368
rect 505590 435334 505642 435368
rect 504962 435278 505642 435334
rect 504962 435244 505016 435278
rect 505050 435244 505106 435278
rect 505140 435244 505196 435278
rect 505230 435244 505286 435278
rect 505320 435244 505376 435278
rect 505410 435244 505466 435278
rect 505500 435244 505556 435278
rect 505590 435244 505642 435278
rect 504962 435188 505642 435244
rect 504962 435154 505016 435188
rect 505050 435154 505106 435188
rect 505140 435154 505196 435188
rect 505230 435154 505286 435188
rect 505320 435154 505376 435188
rect 505410 435154 505466 435188
rect 505500 435154 505556 435188
rect 505590 435154 505642 435188
rect 504962 435098 505642 435154
rect 504962 435064 505016 435098
rect 505050 435064 505106 435098
rect 505140 435064 505196 435098
rect 505230 435064 505286 435098
rect 505320 435064 505376 435098
rect 505410 435064 505466 435098
rect 505500 435064 505556 435098
rect 505590 435064 505642 435098
rect 504962 435008 505642 435064
rect 504962 434974 505016 435008
rect 505050 434974 505106 435008
rect 505140 434974 505196 435008
rect 505230 434974 505286 435008
rect 505320 434974 505376 435008
rect 505410 434974 505466 435008
rect 505500 434974 505556 435008
rect 505590 434974 505642 435008
rect 504962 434922 505642 434974
rect 506250 435548 506930 435602
rect 506250 435514 506304 435548
rect 506338 435514 506394 435548
rect 506428 435514 506484 435548
rect 506518 435514 506574 435548
rect 506608 435514 506664 435548
rect 506698 435514 506754 435548
rect 506788 435514 506844 435548
rect 506878 435514 506930 435548
rect 506250 435458 506930 435514
rect 506250 435424 506304 435458
rect 506338 435424 506394 435458
rect 506428 435424 506484 435458
rect 506518 435424 506574 435458
rect 506608 435424 506664 435458
rect 506698 435424 506754 435458
rect 506788 435424 506844 435458
rect 506878 435424 506930 435458
rect 506250 435368 506930 435424
rect 506250 435334 506304 435368
rect 506338 435334 506394 435368
rect 506428 435334 506484 435368
rect 506518 435334 506574 435368
rect 506608 435334 506664 435368
rect 506698 435334 506754 435368
rect 506788 435334 506844 435368
rect 506878 435334 506930 435368
rect 506250 435278 506930 435334
rect 506250 435244 506304 435278
rect 506338 435244 506394 435278
rect 506428 435244 506484 435278
rect 506518 435244 506574 435278
rect 506608 435244 506664 435278
rect 506698 435244 506754 435278
rect 506788 435244 506844 435278
rect 506878 435244 506930 435278
rect 506250 435188 506930 435244
rect 506250 435154 506304 435188
rect 506338 435154 506394 435188
rect 506428 435154 506484 435188
rect 506518 435154 506574 435188
rect 506608 435154 506664 435188
rect 506698 435154 506754 435188
rect 506788 435154 506844 435188
rect 506878 435154 506930 435188
rect 506250 435098 506930 435154
rect 506250 435064 506304 435098
rect 506338 435064 506394 435098
rect 506428 435064 506484 435098
rect 506518 435064 506574 435098
rect 506608 435064 506664 435098
rect 506698 435064 506754 435098
rect 506788 435064 506844 435098
rect 506878 435064 506930 435098
rect 506250 435008 506930 435064
rect 506250 434974 506304 435008
rect 506338 434974 506394 435008
rect 506428 434974 506484 435008
rect 506518 434974 506574 435008
rect 506608 434974 506664 435008
rect 506698 434974 506754 435008
rect 506788 434974 506844 435008
rect 506878 434974 506930 435008
rect 506250 434922 506930 434974
rect 507538 435548 508218 435602
rect 507538 435514 507592 435548
rect 507626 435514 507682 435548
rect 507716 435514 507772 435548
rect 507806 435514 507862 435548
rect 507896 435514 507952 435548
rect 507986 435514 508042 435548
rect 508076 435514 508132 435548
rect 508166 435514 508218 435548
rect 507538 435458 508218 435514
rect 507538 435424 507592 435458
rect 507626 435424 507682 435458
rect 507716 435424 507772 435458
rect 507806 435424 507862 435458
rect 507896 435424 507952 435458
rect 507986 435424 508042 435458
rect 508076 435424 508132 435458
rect 508166 435424 508218 435458
rect 507538 435368 508218 435424
rect 507538 435334 507592 435368
rect 507626 435334 507682 435368
rect 507716 435334 507772 435368
rect 507806 435334 507862 435368
rect 507896 435334 507952 435368
rect 507986 435334 508042 435368
rect 508076 435334 508132 435368
rect 508166 435334 508218 435368
rect 507538 435278 508218 435334
rect 507538 435244 507592 435278
rect 507626 435244 507682 435278
rect 507716 435244 507772 435278
rect 507806 435244 507862 435278
rect 507896 435244 507952 435278
rect 507986 435244 508042 435278
rect 508076 435244 508132 435278
rect 508166 435244 508218 435278
rect 507538 435188 508218 435244
rect 507538 435154 507592 435188
rect 507626 435154 507682 435188
rect 507716 435154 507772 435188
rect 507806 435154 507862 435188
rect 507896 435154 507952 435188
rect 507986 435154 508042 435188
rect 508076 435154 508132 435188
rect 508166 435154 508218 435188
rect 507538 435098 508218 435154
rect 507538 435064 507592 435098
rect 507626 435064 507682 435098
rect 507716 435064 507772 435098
rect 507806 435064 507862 435098
rect 507896 435064 507952 435098
rect 507986 435064 508042 435098
rect 508076 435064 508132 435098
rect 508166 435064 508218 435098
rect 507538 435008 508218 435064
rect 507538 434974 507592 435008
rect 507626 434974 507682 435008
rect 507716 434974 507772 435008
rect 507806 434974 507862 435008
rect 507896 434974 507952 435008
rect 507986 434974 508042 435008
rect 508076 434974 508132 435008
rect 508166 434974 508218 435008
rect 507538 434922 508218 434974
rect 508826 435548 509506 435602
rect 508826 435514 508880 435548
rect 508914 435514 508970 435548
rect 509004 435514 509060 435548
rect 509094 435514 509150 435548
rect 509184 435514 509240 435548
rect 509274 435514 509330 435548
rect 509364 435514 509420 435548
rect 509454 435514 509506 435548
rect 508826 435458 509506 435514
rect 508826 435424 508880 435458
rect 508914 435424 508970 435458
rect 509004 435424 509060 435458
rect 509094 435424 509150 435458
rect 509184 435424 509240 435458
rect 509274 435424 509330 435458
rect 509364 435424 509420 435458
rect 509454 435424 509506 435458
rect 508826 435368 509506 435424
rect 508826 435334 508880 435368
rect 508914 435334 508970 435368
rect 509004 435334 509060 435368
rect 509094 435334 509150 435368
rect 509184 435334 509240 435368
rect 509274 435334 509330 435368
rect 509364 435334 509420 435368
rect 509454 435334 509506 435368
rect 508826 435278 509506 435334
rect 508826 435244 508880 435278
rect 508914 435244 508970 435278
rect 509004 435244 509060 435278
rect 509094 435244 509150 435278
rect 509184 435244 509240 435278
rect 509274 435244 509330 435278
rect 509364 435244 509420 435278
rect 509454 435244 509506 435278
rect 508826 435188 509506 435244
rect 508826 435154 508880 435188
rect 508914 435154 508970 435188
rect 509004 435154 509060 435188
rect 509094 435154 509150 435188
rect 509184 435154 509240 435188
rect 509274 435154 509330 435188
rect 509364 435154 509420 435188
rect 509454 435154 509506 435188
rect 508826 435098 509506 435154
rect 508826 435064 508880 435098
rect 508914 435064 508970 435098
rect 509004 435064 509060 435098
rect 509094 435064 509150 435098
rect 509184 435064 509240 435098
rect 509274 435064 509330 435098
rect 509364 435064 509420 435098
rect 509454 435064 509506 435098
rect 508826 435008 509506 435064
rect 508826 434974 508880 435008
rect 508914 434974 508970 435008
rect 509004 434974 509060 435008
rect 509094 434974 509150 435008
rect 509184 434974 509240 435008
rect 509274 434974 509330 435008
rect 509364 434974 509420 435008
rect 509454 434974 509506 435008
rect 508826 434922 509506 434974
rect 510114 435548 510794 435602
rect 510114 435514 510168 435548
rect 510202 435514 510258 435548
rect 510292 435514 510348 435548
rect 510382 435514 510438 435548
rect 510472 435514 510528 435548
rect 510562 435514 510618 435548
rect 510652 435514 510708 435548
rect 510742 435514 510794 435548
rect 510114 435458 510794 435514
rect 510114 435424 510168 435458
rect 510202 435424 510258 435458
rect 510292 435424 510348 435458
rect 510382 435424 510438 435458
rect 510472 435424 510528 435458
rect 510562 435424 510618 435458
rect 510652 435424 510708 435458
rect 510742 435424 510794 435458
rect 510114 435368 510794 435424
rect 510114 435334 510168 435368
rect 510202 435334 510258 435368
rect 510292 435334 510348 435368
rect 510382 435334 510438 435368
rect 510472 435334 510528 435368
rect 510562 435334 510618 435368
rect 510652 435334 510708 435368
rect 510742 435334 510794 435368
rect 510114 435278 510794 435334
rect 510114 435244 510168 435278
rect 510202 435244 510258 435278
rect 510292 435244 510348 435278
rect 510382 435244 510438 435278
rect 510472 435244 510528 435278
rect 510562 435244 510618 435278
rect 510652 435244 510708 435278
rect 510742 435244 510794 435278
rect 510114 435188 510794 435244
rect 510114 435154 510168 435188
rect 510202 435154 510258 435188
rect 510292 435154 510348 435188
rect 510382 435154 510438 435188
rect 510472 435154 510528 435188
rect 510562 435154 510618 435188
rect 510652 435154 510708 435188
rect 510742 435154 510794 435188
rect 510114 435098 510794 435154
rect 510114 435064 510168 435098
rect 510202 435064 510258 435098
rect 510292 435064 510348 435098
rect 510382 435064 510438 435098
rect 510472 435064 510528 435098
rect 510562 435064 510618 435098
rect 510652 435064 510708 435098
rect 510742 435064 510794 435098
rect 510114 435008 510794 435064
rect 510114 434974 510168 435008
rect 510202 434974 510258 435008
rect 510292 434974 510348 435008
rect 510382 434974 510438 435008
rect 510472 434974 510528 435008
rect 510562 434974 510618 435008
rect 510652 434974 510708 435008
rect 510742 434974 510794 435008
rect 510114 434922 510794 434974
rect 511402 435548 512082 435602
rect 511402 435514 511456 435548
rect 511490 435514 511546 435548
rect 511580 435514 511636 435548
rect 511670 435514 511726 435548
rect 511760 435514 511816 435548
rect 511850 435514 511906 435548
rect 511940 435514 511996 435548
rect 512030 435514 512082 435548
rect 511402 435458 512082 435514
rect 511402 435424 511456 435458
rect 511490 435424 511546 435458
rect 511580 435424 511636 435458
rect 511670 435424 511726 435458
rect 511760 435424 511816 435458
rect 511850 435424 511906 435458
rect 511940 435424 511996 435458
rect 512030 435424 512082 435458
rect 511402 435368 512082 435424
rect 511402 435334 511456 435368
rect 511490 435334 511546 435368
rect 511580 435334 511636 435368
rect 511670 435334 511726 435368
rect 511760 435334 511816 435368
rect 511850 435334 511906 435368
rect 511940 435334 511996 435368
rect 512030 435334 512082 435368
rect 511402 435278 512082 435334
rect 511402 435244 511456 435278
rect 511490 435244 511546 435278
rect 511580 435244 511636 435278
rect 511670 435244 511726 435278
rect 511760 435244 511816 435278
rect 511850 435244 511906 435278
rect 511940 435244 511996 435278
rect 512030 435244 512082 435278
rect 511402 435188 512082 435244
rect 511402 435154 511456 435188
rect 511490 435154 511546 435188
rect 511580 435154 511636 435188
rect 511670 435154 511726 435188
rect 511760 435154 511816 435188
rect 511850 435154 511906 435188
rect 511940 435154 511996 435188
rect 512030 435154 512082 435188
rect 511402 435098 512082 435154
rect 511402 435064 511456 435098
rect 511490 435064 511546 435098
rect 511580 435064 511636 435098
rect 511670 435064 511726 435098
rect 511760 435064 511816 435098
rect 511850 435064 511906 435098
rect 511940 435064 511996 435098
rect 512030 435064 512082 435098
rect 511402 435008 512082 435064
rect 511402 434974 511456 435008
rect 511490 434974 511546 435008
rect 511580 434974 511636 435008
rect 511670 434974 511726 435008
rect 511760 434974 511816 435008
rect 511850 434974 511906 435008
rect 511940 434974 511996 435008
rect 512030 434974 512082 435008
rect 511402 434922 512082 434974
rect 512690 435548 513370 435602
rect 512690 435514 512744 435548
rect 512778 435514 512834 435548
rect 512868 435514 512924 435548
rect 512958 435514 513014 435548
rect 513048 435514 513104 435548
rect 513138 435514 513194 435548
rect 513228 435514 513284 435548
rect 513318 435514 513370 435548
rect 512690 435458 513370 435514
rect 512690 435424 512744 435458
rect 512778 435424 512834 435458
rect 512868 435424 512924 435458
rect 512958 435424 513014 435458
rect 513048 435424 513104 435458
rect 513138 435424 513194 435458
rect 513228 435424 513284 435458
rect 513318 435424 513370 435458
rect 512690 435368 513370 435424
rect 512690 435334 512744 435368
rect 512778 435334 512834 435368
rect 512868 435334 512924 435368
rect 512958 435334 513014 435368
rect 513048 435334 513104 435368
rect 513138 435334 513194 435368
rect 513228 435334 513284 435368
rect 513318 435334 513370 435368
rect 512690 435278 513370 435334
rect 512690 435244 512744 435278
rect 512778 435244 512834 435278
rect 512868 435244 512924 435278
rect 512958 435244 513014 435278
rect 513048 435244 513104 435278
rect 513138 435244 513194 435278
rect 513228 435244 513284 435278
rect 513318 435244 513370 435278
rect 512690 435188 513370 435244
rect 512690 435154 512744 435188
rect 512778 435154 512834 435188
rect 512868 435154 512924 435188
rect 512958 435154 513014 435188
rect 513048 435154 513104 435188
rect 513138 435154 513194 435188
rect 513228 435154 513284 435188
rect 513318 435154 513370 435188
rect 512690 435098 513370 435154
rect 512690 435064 512744 435098
rect 512778 435064 512834 435098
rect 512868 435064 512924 435098
rect 512958 435064 513014 435098
rect 513048 435064 513104 435098
rect 513138 435064 513194 435098
rect 513228 435064 513284 435098
rect 513318 435064 513370 435098
rect 512690 435008 513370 435064
rect 512690 434974 512744 435008
rect 512778 434974 512834 435008
rect 512868 434974 512924 435008
rect 512958 434974 513014 435008
rect 513048 434974 513104 435008
rect 513138 434974 513194 435008
rect 513228 434974 513284 435008
rect 513318 434974 513370 435008
rect 512690 434922 513370 434974
rect 503674 434260 504354 434314
rect 503674 434226 503728 434260
rect 503762 434226 503818 434260
rect 503852 434226 503908 434260
rect 503942 434226 503998 434260
rect 504032 434226 504088 434260
rect 504122 434226 504178 434260
rect 504212 434226 504268 434260
rect 504302 434226 504354 434260
rect 503674 434170 504354 434226
rect 503674 434136 503728 434170
rect 503762 434136 503818 434170
rect 503852 434136 503908 434170
rect 503942 434136 503998 434170
rect 504032 434136 504088 434170
rect 504122 434136 504178 434170
rect 504212 434136 504268 434170
rect 504302 434136 504354 434170
rect 503674 434080 504354 434136
rect 503674 434046 503728 434080
rect 503762 434046 503818 434080
rect 503852 434046 503908 434080
rect 503942 434046 503998 434080
rect 504032 434046 504088 434080
rect 504122 434046 504178 434080
rect 504212 434046 504268 434080
rect 504302 434046 504354 434080
rect 503674 433990 504354 434046
rect 503674 433956 503728 433990
rect 503762 433956 503818 433990
rect 503852 433956 503908 433990
rect 503942 433956 503998 433990
rect 504032 433956 504088 433990
rect 504122 433956 504178 433990
rect 504212 433956 504268 433990
rect 504302 433956 504354 433990
rect 503674 433900 504354 433956
rect 503674 433866 503728 433900
rect 503762 433866 503818 433900
rect 503852 433866 503908 433900
rect 503942 433866 503998 433900
rect 504032 433866 504088 433900
rect 504122 433866 504178 433900
rect 504212 433866 504268 433900
rect 504302 433866 504354 433900
rect 503674 433810 504354 433866
rect 503674 433776 503728 433810
rect 503762 433776 503818 433810
rect 503852 433776 503908 433810
rect 503942 433776 503998 433810
rect 504032 433776 504088 433810
rect 504122 433776 504178 433810
rect 504212 433776 504268 433810
rect 504302 433776 504354 433810
rect 503674 433720 504354 433776
rect 503674 433686 503728 433720
rect 503762 433686 503818 433720
rect 503852 433686 503908 433720
rect 503942 433686 503998 433720
rect 504032 433686 504088 433720
rect 504122 433686 504178 433720
rect 504212 433686 504268 433720
rect 504302 433686 504354 433720
rect 503674 433634 504354 433686
rect 504962 434260 505642 434314
rect 504962 434226 505016 434260
rect 505050 434226 505106 434260
rect 505140 434226 505196 434260
rect 505230 434226 505286 434260
rect 505320 434226 505376 434260
rect 505410 434226 505466 434260
rect 505500 434226 505556 434260
rect 505590 434226 505642 434260
rect 504962 434170 505642 434226
rect 504962 434136 505016 434170
rect 505050 434136 505106 434170
rect 505140 434136 505196 434170
rect 505230 434136 505286 434170
rect 505320 434136 505376 434170
rect 505410 434136 505466 434170
rect 505500 434136 505556 434170
rect 505590 434136 505642 434170
rect 504962 434080 505642 434136
rect 504962 434046 505016 434080
rect 505050 434046 505106 434080
rect 505140 434046 505196 434080
rect 505230 434046 505286 434080
rect 505320 434046 505376 434080
rect 505410 434046 505466 434080
rect 505500 434046 505556 434080
rect 505590 434046 505642 434080
rect 504962 433990 505642 434046
rect 504962 433956 505016 433990
rect 505050 433956 505106 433990
rect 505140 433956 505196 433990
rect 505230 433956 505286 433990
rect 505320 433956 505376 433990
rect 505410 433956 505466 433990
rect 505500 433956 505556 433990
rect 505590 433956 505642 433990
rect 504962 433900 505642 433956
rect 504962 433866 505016 433900
rect 505050 433866 505106 433900
rect 505140 433866 505196 433900
rect 505230 433866 505286 433900
rect 505320 433866 505376 433900
rect 505410 433866 505466 433900
rect 505500 433866 505556 433900
rect 505590 433866 505642 433900
rect 504962 433810 505642 433866
rect 504962 433776 505016 433810
rect 505050 433776 505106 433810
rect 505140 433776 505196 433810
rect 505230 433776 505286 433810
rect 505320 433776 505376 433810
rect 505410 433776 505466 433810
rect 505500 433776 505556 433810
rect 505590 433776 505642 433810
rect 504962 433720 505642 433776
rect 504962 433686 505016 433720
rect 505050 433686 505106 433720
rect 505140 433686 505196 433720
rect 505230 433686 505286 433720
rect 505320 433686 505376 433720
rect 505410 433686 505466 433720
rect 505500 433686 505556 433720
rect 505590 433686 505642 433720
rect 504962 433634 505642 433686
rect 506250 434260 506930 434314
rect 506250 434226 506304 434260
rect 506338 434226 506394 434260
rect 506428 434226 506484 434260
rect 506518 434226 506574 434260
rect 506608 434226 506664 434260
rect 506698 434226 506754 434260
rect 506788 434226 506844 434260
rect 506878 434226 506930 434260
rect 506250 434170 506930 434226
rect 506250 434136 506304 434170
rect 506338 434136 506394 434170
rect 506428 434136 506484 434170
rect 506518 434136 506574 434170
rect 506608 434136 506664 434170
rect 506698 434136 506754 434170
rect 506788 434136 506844 434170
rect 506878 434136 506930 434170
rect 506250 434080 506930 434136
rect 506250 434046 506304 434080
rect 506338 434046 506394 434080
rect 506428 434046 506484 434080
rect 506518 434046 506574 434080
rect 506608 434046 506664 434080
rect 506698 434046 506754 434080
rect 506788 434046 506844 434080
rect 506878 434046 506930 434080
rect 506250 433990 506930 434046
rect 506250 433956 506304 433990
rect 506338 433956 506394 433990
rect 506428 433956 506484 433990
rect 506518 433956 506574 433990
rect 506608 433956 506664 433990
rect 506698 433956 506754 433990
rect 506788 433956 506844 433990
rect 506878 433956 506930 433990
rect 506250 433900 506930 433956
rect 506250 433866 506304 433900
rect 506338 433866 506394 433900
rect 506428 433866 506484 433900
rect 506518 433866 506574 433900
rect 506608 433866 506664 433900
rect 506698 433866 506754 433900
rect 506788 433866 506844 433900
rect 506878 433866 506930 433900
rect 506250 433810 506930 433866
rect 506250 433776 506304 433810
rect 506338 433776 506394 433810
rect 506428 433776 506484 433810
rect 506518 433776 506574 433810
rect 506608 433776 506664 433810
rect 506698 433776 506754 433810
rect 506788 433776 506844 433810
rect 506878 433776 506930 433810
rect 506250 433720 506930 433776
rect 506250 433686 506304 433720
rect 506338 433686 506394 433720
rect 506428 433686 506484 433720
rect 506518 433686 506574 433720
rect 506608 433686 506664 433720
rect 506698 433686 506754 433720
rect 506788 433686 506844 433720
rect 506878 433686 506930 433720
rect 506250 433634 506930 433686
rect 507538 434260 508218 434314
rect 507538 434226 507592 434260
rect 507626 434226 507682 434260
rect 507716 434226 507772 434260
rect 507806 434226 507862 434260
rect 507896 434226 507952 434260
rect 507986 434226 508042 434260
rect 508076 434226 508132 434260
rect 508166 434226 508218 434260
rect 507538 434170 508218 434226
rect 507538 434136 507592 434170
rect 507626 434136 507682 434170
rect 507716 434136 507772 434170
rect 507806 434136 507862 434170
rect 507896 434136 507952 434170
rect 507986 434136 508042 434170
rect 508076 434136 508132 434170
rect 508166 434136 508218 434170
rect 507538 434080 508218 434136
rect 507538 434046 507592 434080
rect 507626 434046 507682 434080
rect 507716 434046 507772 434080
rect 507806 434046 507862 434080
rect 507896 434046 507952 434080
rect 507986 434046 508042 434080
rect 508076 434046 508132 434080
rect 508166 434046 508218 434080
rect 507538 433990 508218 434046
rect 507538 433956 507592 433990
rect 507626 433956 507682 433990
rect 507716 433956 507772 433990
rect 507806 433956 507862 433990
rect 507896 433956 507952 433990
rect 507986 433956 508042 433990
rect 508076 433956 508132 433990
rect 508166 433956 508218 433990
rect 507538 433900 508218 433956
rect 507538 433866 507592 433900
rect 507626 433866 507682 433900
rect 507716 433866 507772 433900
rect 507806 433866 507862 433900
rect 507896 433866 507952 433900
rect 507986 433866 508042 433900
rect 508076 433866 508132 433900
rect 508166 433866 508218 433900
rect 507538 433810 508218 433866
rect 507538 433776 507592 433810
rect 507626 433776 507682 433810
rect 507716 433776 507772 433810
rect 507806 433776 507862 433810
rect 507896 433776 507952 433810
rect 507986 433776 508042 433810
rect 508076 433776 508132 433810
rect 508166 433776 508218 433810
rect 507538 433720 508218 433776
rect 507538 433686 507592 433720
rect 507626 433686 507682 433720
rect 507716 433686 507772 433720
rect 507806 433686 507862 433720
rect 507896 433686 507952 433720
rect 507986 433686 508042 433720
rect 508076 433686 508132 433720
rect 508166 433686 508218 433720
rect 507538 433634 508218 433686
rect 508826 434260 509506 434314
rect 508826 434226 508880 434260
rect 508914 434226 508970 434260
rect 509004 434226 509060 434260
rect 509094 434226 509150 434260
rect 509184 434226 509240 434260
rect 509274 434226 509330 434260
rect 509364 434226 509420 434260
rect 509454 434226 509506 434260
rect 508826 434170 509506 434226
rect 508826 434136 508880 434170
rect 508914 434136 508970 434170
rect 509004 434136 509060 434170
rect 509094 434136 509150 434170
rect 509184 434136 509240 434170
rect 509274 434136 509330 434170
rect 509364 434136 509420 434170
rect 509454 434136 509506 434170
rect 508826 434080 509506 434136
rect 508826 434046 508880 434080
rect 508914 434046 508970 434080
rect 509004 434046 509060 434080
rect 509094 434046 509150 434080
rect 509184 434046 509240 434080
rect 509274 434046 509330 434080
rect 509364 434046 509420 434080
rect 509454 434046 509506 434080
rect 508826 433990 509506 434046
rect 508826 433956 508880 433990
rect 508914 433956 508970 433990
rect 509004 433956 509060 433990
rect 509094 433956 509150 433990
rect 509184 433956 509240 433990
rect 509274 433956 509330 433990
rect 509364 433956 509420 433990
rect 509454 433956 509506 433990
rect 508826 433900 509506 433956
rect 508826 433866 508880 433900
rect 508914 433866 508970 433900
rect 509004 433866 509060 433900
rect 509094 433866 509150 433900
rect 509184 433866 509240 433900
rect 509274 433866 509330 433900
rect 509364 433866 509420 433900
rect 509454 433866 509506 433900
rect 508826 433810 509506 433866
rect 508826 433776 508880 433810
rect 508914 433776 508970 433810
rect 509004 433776 509060 433810
rect 509094 433776 509150 433810
rect 509184 433776 509240 433810
rect 509274 433776 509330 433810
rect 509364 433776 509420 433810
rect 509454 433776 509506 433810
rect 508826 433720 509506 433776
rect 508826 433686 508880 433720
rect 508914 433686 508970 433720
rect 509004 433686 509060 433720
rect 509094 433686 509150 433720
rect 509184 433686 509240 433720
rect 509274 433686 509330 433720
rect 509364 433686 509420 433720
rect 509454 433686 509506 433720
rect 508826 433634 509506 433686
rect 510114 434260 510794 434314
rect 510114 434226 510168 434260
rect 510202 434226 510258 434260
rect 510292 434226 510348 434260
rect 510382 434226 510438 434260
rect 510472 434226 510528 434260
rect 510562 434226 510618 434260
rect 510652 434226 510708 434260
rect 510742 434226 510794 434260
rect 510114 434170 510794 434226
rect 510114 434136 510168 434170
rect 510202 434136 510258 434170
rect 510292 434136 510348 434170
rect 510382 434136 510438 434170
rect 510472 434136 510528 434170
rect 510562 434136 510618 434170
rect 510652 434136 510708 434170
rect 510742 434136 510794 434170
rect 510114 434080 510794 434136
rect 510114 434046 510168 434080
rect 510202 434046 510258 434080
rect 510292 434046 510348 434080
rect 510382 434046 510438 434080
rect 510472 434046 510528 434080
rect 510562 434046 510618 434080
rect 510652 434046 510708 434080
rect 510742 434046 510794 434080
rect 510114 433990 510794 434046
rect 510114 433956 510168 433990
rect 510202 433956 510258 433990
rect 510292 433956 510348 433990
rect 510382 433956 510438 433990
rect 510472 433956 510528 433990
rect 510562 433956 510618 433990
rect 510652 433956 510708 433990
rect 510742 433956 510794 433990
rect 510114 433900 510794 433956
rect 510114 433866 510168 433900
rect 510202 433866 510258 433900
rect 510292 433866 510348 433900
rect 510382 433866 510438 433900
rect 510472 433866 510528 433900
rect 510562 433866 510618 433900
rect 510652 433866 510708 433900
rect 510742 433866 510794 433900
rect 510114 433810 510794 433866
rect 510114 433776 510168 433810
rect 510202 433776 510258 433810
rect 510292 433776 510348 433810
rect 510382 433776 510438 433810
rect 510472 433776 510528 433810
rect 510562 433776 510618 433810
rect 510652 433776 510708 433810
rect 510742 433776 510794 433810
rect 510114 433720 510794 433776
rect 510114 433686 510168 433720
rect 510202 433686 510258 433720
rect 510292 433686 510348 433720
rect 510382 433686 510438 433720
rect 510472 433686 510528 433720
rect 510562 433686 510618 433720
rect 510652 433686 510708 433720
rect 510742 433686 510794 433720
rect 510114 433634 510794 433686
rect 511402 434260 512082 434314
rect 511402 434226 511456 434260
rect 511490 434226 511546 434260
rect 511580 434226 511636 434260
rect 511670 434226 511726 434260
rect 511760 434226 511816 434260
rect 511850 434226 511906 434260
rect 511940 434226 511996 434260
rect 512030 434226 512082 434260
rect 511402 434170 512082 434226
rect 511402 434136 511456 434170
rect 511490 434136 511546 434170
rect 511580 434136 511636 434170
rect 511670 434136 511726 434170
rect 511760 434136 511816 434170
rect 511850 434136 511906 434170
rect 511940 434136 511996 434170
rect 512030 434136 512082 434170
rect 511402 434080 512082 434136
rect 511402 434046 511456 434080
rect 511490 434046 511546 434080
rect 511580 434046 511636 434080
rect 511670 434046 511726 434080
rect 511760 434046 511816 434080
rect 511850 434046 511906 434080
rect 511940 434046 511996 434080
rect 512030 434046 512082 434080
rect 511402 433990 512082 434046
rect 511402 433956 511456 433990
rect 511490 433956 511546 433990
rect 511580 433956 511636 433990
rect 511670 433956 511726 433990
rect 511760 433956 511816 433990
rect 511850 433956 511906 433990
rect 511940 433956 511996 433990
rect 512030 433956 512082 433990
rect 511402 433900 512082 433956
rect 511402 433866 511456 433900
rect 511490 433866 511546 433900
rect 511580 433866 511636 433900
rect 511670 433866 511726 433900
rect 511760 433866 511816 433900
rect 511850 433866 511906 433900
rect 511940 433866 511996 433900
rect 512030 433866 512082 433900
rect 511402 433810 512082 433866
rect 511402 433776 511456 433810
rect 511490 433776 511546 433810
rect 511580 433776 511636 433810
rect 511670 433776 511726 433810
rect 511760 433776 511816 433810
rect 511850 433776 511906 433810
rect 511940 433776 511996 433810
rect 512030 433776 512082 433810
rect 511402 433720 512082 433776
rect 511402 433686 511456 433720
rect 511490 433686 511546 433720
rect 511580 433686 511636 433720
rect 511670 433686 511726 433720
rect 511760 433686 511816 433720
rect 511850 433686 511906 433720
rect 511940 433686 511996 433720
rect 512030 433686 512082 433720
rect 511402 433634 512082 433686
rect 512690 434260 513370 434314
rect 512690 434226 512744 434260
rect 512778 434226 512834 434260
rect 512868 434226 512924 434260
rect 512958 434226 513014 434260
rect 513048 434226 513104 434260
rect 513138 434226 513194 434260
rect 513228 434226 513284 434260
rect 513318 434226 513370 434260
rect 512690 434170 513370 434226
rect 512690 434136 512744 434170
rect 512778 434136 512834 434170
rect 512868 434136 512924 434170
rect 512958 434136 513014 434170
rect 513048 434136 513104 434170
rect 513138 434136 513194 434170
rect 513228 434136 513284 434170
rect 513318 434136 513370 434170
rect 512690 434080 513370 434136
rect 512690 434046 512744 434080
rect 512778 434046 512834 434080
rect 512868 434046 512924 434080
rect 512958 434046 513014 434080
rect 513048 434046 513104 434080
rect 513138 434046 513194 434080
rect 513228 434046 513284 434080
rect 513318 434046 513370 434080
rect 512690 433990 513370 434046
rect 512690 433956 512744 433990
rect 512778 433956 512834 433990
rect 512868 433956 512924 433990
rect 512958 433956 513014 433990
rect 513048 433956 513104 433990
rect 513138 433956 513194 433990
rect 513228 433956 513284 433990
rect 513318 433956 513370 433990
rect 512690 433900 513370 433956
rect 512690 433866 512744 433900
rect 512778 433866 512834 433900
rect 512868 433866 512924 433900
rect 512958 433866 513014 433900
rect 513048 433866 513104 433900
rect 513138 433866 513194 433900
rect 513228 433866 513284 433900
rect 513318 433866 513370 433900
rect 512690 433810 513370 433866
rect 512690 433776 512744 433810
rect 512778 433776 512834 433810
rect 512868 433776 512924 433810
rect 512958 433776 513014 433810
rect 513048 433776 513104 433810
rect 513138 433776 513194 433810
rect 513228 433776 513284 433810
rect 513318 433776 513370 433810
rect 512690 433720 513370 433776
rect 512690 433686 512744 433720
rect 512778 433686 512834 433720
rect 512868 433686 512924 433720
rect 512958 433686 513014 433720
rect 513048 433686 513104 433720
rect 513138 433686 513194 433720
rect 513228 433686 513284 433720
rect 513318 433686 513370 433720
rect 512690 433634 513370 433686
rect 503674 432972 504354 433026
rect 503674 432938 503728 432972
rect 503762 432938 503818 432972
rect 503852 432938 503908 432972
rect 503942 432938 503998 432972
rect 504032 432938 504088 432972
rect 504122 432938 504178 432972
rect 504212 432938 504268 432972
rect 504302 432938 504354 432972
rect 503674 432882 504354 432938
rect 503674 432848 503728 432882
rect 503762 432848 503818 432882
rect 503852 432848 503908 432882
rect 503942 432848 503998 432882
rect 504032 432848 504088 432882
rect 504122 432848 504178 432882
rect 504212 432848 504268 432882
rect 504302 432848 504354 432882
rect 503674 432792 504354 432848
rect 503674 432758 503728 432792
rect 503762 432758 503818 432792
rect 503852 432758 503908 432792
rect 503942 432758 503998 432792
rect 504032 432758 504088 432792
rect 504122 432758 504178 432792
rect 504212 432758 504268 432792
rect 504302 432758 504354 432792
rect 503674 432702 504354 432758
rect 503674 432668 503728 432702
rect 503762 432668 503818 432702
rect 503852 432668 503908 432702
rect 503942 432668 503998 432702
rect 504032 432668 504088 432702
rect 504122 432668 504178 432702
rect 504212 432668 504268 432702
rect 504302 432668 504354 432702
rect 503674 432612 504354 432668
rect 503674 432578 503728 432612
rect 503762 432578 503818 432612
rect 503852 432578 503908 432612
rect 503942 432578 503998 432612
rect 504032 432578 504088 432612
rect 504122 432578 504178 432612
rect 504212 432578 504268 432612
rect 504302 432578 504354 432612
rect 503674 432522 504354 432578
rect 503674 432488 503728 432522
rect 503762 432488 503818 432522
rect 503852 432488 503908 432522
rect 503942 432488 503998 432522
rect 504032 432488 504088 432522
rect 504122 432488 504178 432522
rect 504212 432488 504268 432522
rect 504302 432488 504354 432522
rect 503674 432432 504354 432488
rect 503674 432398 503728 432432
rect 503762 432398 503818 432432
rect 503852 432398 503908 432432
rect 503942 432398 503998 432432
rect 504032 432398 504088 432432
rect 504122 432398 504178 432432
rect 504212 432398 504268 432432
rect 504302 432398 504354 432432
rect 503674 432346 504354 432398
rect 504962 432972 505642 433026
rect 504962 432938 505016 432972
rect 505050 432938 505106 432972
rect 505140 432938 505196 432972
rect 505230 432938 505286 432972
rect 505320 432938 505376 432972
rect 505410 432938 505466 432972
rect 505500 432938 505556 432972
rect 505590 432938 505642 432972
rect 504962 432882 505642 432938
rect 504962 432848 505016 432882
rect 505050 432848 505106 432882
rect 505140 432848 505196 432882
rect 505230 432848 505286 432882
rect 505320 432848 505376 432882
rect 505410 432848 505466 432882
rect 505500 432848 505556 432882
rect 505590 432848 505642 432882
rect 504962 432792 505642 432848
rect 504962 432758 505016 432792
rect 505050 432758 505106 432792
rect 505140 432758 505196 432792
rect 505230 432758 505286 432792
rect 505320 432758 505376 432792
rect 505410 432758 505466 432792
rect 505500 432758 505556 432792
rect 505590 432758 505642 432792
rect 504962 432702 505642 432758
rect 504962 432668 505016 432702
rect 505050 432668 505106 432702
rect 505140 432668 505196 432702
rect 505230 432668 505286 432702
rect 505320 432668 505376 432702
rect 505410 432668 505466 432702
rect 505500 432668 505556 432702
rect 505590 432668 505642 432702
rect 504962 432612 505642 432668
rect 504962 432578 505016 432612
rect 505050 432578 505106 432612
rect 505140 432578 505196 432612
rect 505230 432578 505286 432612
rect 505320 432578 505376 432612
rect 505410 432578 505466 432612
rect 505500 432578 505556 432612
rect 505590 432578 505642 432612
rect 504962 432522 505642 432578
rect 504962 432488 505016 432522
rect 505050 432488 505106 432522
rect 505140 432488 505196 432522
rect 505230 432488 505286 432522
rect 505320 432488 505376 432522
rect 505410 432488 505466 432522
rect 505500 432488 505556 432522
rect 505590 432488 505642 432522
rect 504962 432432 505642 432488
rect 504962 432398 505016 432432
rect 505050 432398 505106 432432
rect 505140 432398 505196 432432
rect 505230 432398 505286 432432
rect 505320 432398 505376 432432
rect 505410 432398 505466 432432
rect 505500 432398 505556 432432
rect 505590 432398 505642 432432
rect 504962 432346 505642 432398
rect 506250 432972 506930 433026
rect 506250 432938 506304 432972
rect 506338 432938 506394 432972
rect 506428 432938 506484 432972
rect 506518 432938 506574 432972
rect 506608 432938 506664 432972
rect 506698 432938 506754 432972
rect 506788 432938 506844 432972
rect 506878 432938 506930 432972
rect 506250 432882 506930 432938
rect 506250 432848 506304 432882
rect 506338 432848 506394 432882
rect 506428 432848 506484 432882
rect 506518 432848 506574 432882
rect 506608 432848 506664 432882
rect 506698 432848 506754 432882
rect 506788 432848 506844 432882
rect 506878 432848 506930 432882
rect 506250 432792 506930 432848
rect 506250 432758 506304 432792
rect 506338 432758 506394 432792
rect 506428 432758 506484 432792
rect 506518 432758 506574 432792
rect 506608 432758 506664 432792
rect 506698 432758 506754 432792
rect 506788 432758 506844 432792
rect 506878 432758 506930 432792
rect 506250 432702 506930 432758
rect 506250 432668 506304 432702
rect 506338 432668 506394 432702
rect 506428 432668 506484 432702
rect 506518 432668 506574 432702
rect 506608 432668 506664 432702
rect 506698 432668 506754 432702
rect 506788 432668 506844 432702
rect 506878 432668 506930 432702
rect 506250 432612 506930 432668
rect 506250 432578 506304 432612
rect 506338 432578 506394 432612
rect 506428 432578 506484 432612
rect 506518 432578 506574 432612
rect 506608 432578 506664 432612
rect 506698 432578 506754 432612
rect 506788 432578 506844 432612
rect 506878 432578 506930 432612
rect 506250 432522 506930 432578
rect 506250 432488 506304 432522
rect 506338 432488 506394 432522
rect 506428 432488 506484 432522
rect 506518 432488 506574 432522
rect 506608 432488 506664 432522
rect 506698 432488 506754 432522
rect 506788 432488 506844 432522
rect 506878 432488 506930 432522
rect 506250 432432 506930 432488
rect 506250 432398 506304 432432
rect 506338 432398 506394 432432
rect 506428 432398 506484 432432
rect 506518 432398 506574 432432
rect 506608 432398 506664 432432
rect 506698 432398 506754 432432
rect 506788 432398 506844 432432
rect 506878 432398 506930 432432
rect 506250 432346 506930 432398
rect 507538 432972 508218 433026
rect 507538 432938 507592 432972
rect 507626 432938 507682 432972
rect 507716 432938 507772 432972
rect 507806 432938 507862 432972
rect 507896 432938 507952 432972
rect 507986 432938 508042 432972
rect 508076 432938 508132 432972
rect 508166 432938 508218 432972
rect 507538 432882 508218 432938
rect 507538 432848 507592 432882
rect 507626 432848 507682 432882
rect 507716 432848 507772 432882
rect 507806 432848 507862 432882
rect 507896 432848 507952 432882
rect 507986 432848 508042 432882
rect 508076 432848 508132 432882
rect 508166 432848 508218 432882
rect 507538 432792 508218 432848
rect 507538 432758 507592 432792
rect 507626 432758 507682 432792
rect 507716 432758 507772 432792
rect 507806 432758 507862 432792
rect 507896 432758 507952 432792
rect 507986 432758 508042 432792
rect 508076 432758 508132 432792
rect 508166 432758 508218 432792
rect 507538 432702 508218 432758
rect 507538 432668 507592 432702
rect 507626 432668 507682 432702
rect 507716 432668 507772 432702
rect 507806 432668 507862 432702
rect 507896 432668 507952 432702
rect 507986 432668 508042 432702
rect 508076 432668 508132 432702
rect 508166 432668 508218 432702
rect 507538 432612 508218 432668
rect 507538 432578 507592 432612
rect 507626 432578 507682 432612
rect 507716 432578 507772 432612
rect 507806 432578 507862 432612
rect 507896 432578 507952 432612
rect 507986 432578 508042 432612
rect 508076 432578 508132 432612
rect 508166 432578 508218 432612
rect 507538 432522 508218 432578
rect 507538 432488 507592 432522
rect 507626 432488 507682 432522
rect 507716 432488 507772 432522
rect 507806 432488 507862 432522
rect 507896 432488 507952 432522
rect 507986 432488 508042 432522
rect 508076 432488 508132 432522
rect 508166 432488 508218 432522
rect 507538 432432 508218 432488
rect 507538 432398 507592 432432
rect 507626 432398 507682 432432
rect 507716 432398 507772 432432
rect 507806 432398 507862 432432
rect 507896 432398 507952 432432
rect 507986 432398 508042 432432
rect 508076 432398 508132 432432
rect 508166 432398 508218 432432
rect 507538 432346 508218 432398
rect 508826 432972 509506 433026
rect 508826 432938 508880 432972
rect 508914 432938 508970 432972
rect 509004 432938 509060 432972
rect 509094 432938 509150 432972
rect 509184 432938 509240 432972
rect 509274 432938 509330 432972
rect 509364 432938 509420 432972
rect 509454 432938 509506 432972
rect 508826 432882 509506 432938
rect 508826 432848 508880 432882
rect 508914 432848 508970 432882
rect 509004 432848 509060 432882
rect 509094 432848 509150 432882
rect 509184 432848 509240 432882
rect 509274 432848 509330 432882
rect 509364 432848 509420 432882
rect 509454 432848 509506 432882
rect 508826 432792 509506 432848
rect 508826 432758 508880 432792
rect 508914 432758 508970 432792
rect 509004 432758 509060 432792
rect 509094 432758 509150 432792
rect 509184 432758 509240 432792
rect 509274 432758 509330 432792
rect 509364 432758 509420 432792
rect 509454 432758 509506 432792
rect 508826 432702 509506 432758
rect 508826 432668 508880 432702
rect 508914 432668 508970 432702
rect 509004 432668 509060 432702
rect 509094 432668 509150 432702
rect 509184 432668 509240 432702
rect 509274 432668 509330 432702
rect 509364 432668 509420 432702
rect 509454 432668 509506 432702
rect 508826 432612 509506 432668
rect 508826 432578 508880 432612
rect 508914 432578 508970 432612
rect 509004 432578 509060 432612
rect 509094 432578 509150 432612
rect 509184 432578 509240 432612
rect 509274 432578 509330 432612
rect 509364 432578 509420 432612
rect 509454 432578 509506 432612
rect 508826 432522 509506 432578
rect 508826 432488 508880 432522
rect 508914 432488 508970 432522
rect 509004 432488 509060 432522
rect 509094 432488 509150 432522
rect 509184 432488 509240 432522
rect 509274 432488 509330 432522
rect 509364 432488 509420 432522
rect 509454 432488 509506 432522
rect 508826 432432 509506 432488
rect 508826 432398 508880 432432
rect 508914 432398 508970 432432
rect 509004 432398 509060 432432
rect 509094 432398 509150 432432
rect 509184 432398 509240 432432
rect 509274 432398 509330 432432
rect 509364 432398 509420 432432
rect 509454 432398 509506 432432
rect 508826 432346 509506 432398
rect 510114 432972 510794 433026
rect 510114 432938 510168 432972
rect 510202 432938 510258 432972
rect 510292 432938 510348 432972
rect 510382 432938 510438 432972
rect 510472 432938 510528 432972
rect 510562 432938 510618 432972
rect 510652 432938 510708 432972
rect 510742 432938 510794 432972
rect 510114 432882 510794 432938
rect 510114 432848 510168 432882
rect 510202 432848 510258 432882
rect 510292 432848 510348 432882
rect 510382 432848 510438 432882
rect 510472 432848 510528 432882
rect 510562 432848 510618 432882
rect 510652 432848 510708 432882
rect 510742 432848 510794 432882
rect 510114 432792 510794 432848
rect 510114 432758 510168 432792
rect 510202 432758 510258 432792
rect 510292 432758 510348 432792
rect 510382 432758 510438 432792
rect 510472 432758 510528 432792
rect 510562 432758 510618 432792
rect 510652 432758 510708 432792
rect 510742 432758 510794 432792
rect 510114 432702 510794 432758
rect 510114 432668 510168 432702
rect 510202 432668 510258 432702
rect 510292 432668 510348 432702
rect 510382 432668 510438 432702
rect 510472 432668 510528 432702
rect 510562 432668 510618 432702
rect 510652 432668 510708 432702
rect 510742 432668 510794 432702
rect 510114 432612 510794 432668
rect 510114 432578 510168 432612
rect 510202 432578 510258 432612
rect 510292 432578 510348 432612
rect 510382 432578 510438 432612
rect 510472 432578 510528 432612
rect 510562 432578 510618 432612
rect 510652 432578 510708 432612
rect 510742 432578 510794 432612
rect 510114 432522 510794 432578
rect 510114 432488 510168 432522
rect 510202 432488 510258 432522
rect 510292 432488 510348 432522
rect 510382 432488 510438 432522
rect 510472 432488 510528 432522
rect 510562 432488 510618 432522
rect 510652 432488 510708 432522
rect 510742 432488 510794 432522
rect 510114 432432 510794 432488
rect 510114 432398 510168 432432
rect 510202 432398 510258 432432
rect 510292 432398 510348 432432
rect 510382 432398 510438 432432
rect 510472 432398 510528 432432
rect 510562 432398 510618 432432
rect 510652 432398 510708 432432
rect 510742 432398 510794 432432
rect 510114 432346 510794 432398
rect 511402 432972 512082 433026
rect 511402 432938 511456 432972
rect 511490 432938 511546 432972
rect 511580 432938 511636 432972
rect 511670 432938 511726 432972
rect 511760 432938 511816 432972
rect 511850 432938 511906 432972
rect 511940 432938 511996 432972
rect 512030 432938 512082 432972
rect 511402 432882 512082 432938
rect 511402 432848 511456 432882
rect 511490 432848 511546 432882
rect 511580 432848 511636 432882
rect 511670 432848 511726 432882
rect 511760 432848 511816 432882
rect 511850 432848 511906 432882
rect 511940 432848 511996 432882
rect 512030 432848 512082 432882
rect 511402 432792 512082 432848
rect 511402 432758 511456 432792
rect 511490 432758 511546 432792
rect 511580 432758 511636 432792
rect 511670 432758 511726 432792
rect 511760 432758 511816 432792
rect 511850 432758 511906 432792
rect 511940 432758 511996 432792
rect 512030 432758 512082 432792
rect 511402 432702 512082 432758
rect 511402 432668 511456 432702
rect 511490 432668 511546 432702
rect 511580 432668 511636 432702
rect 511670 432668 511726 432702
rect 511760 432668 511816 432702
rect 511850 432668 511906 432702
rect 511940 432668 511996 432702
rect 512030 432668 512082 432702
rect 511402 432612 512082 432668
rect 511402 432578 511456 432612
rect 511490 432578 511546 432612
rect 511580 432578 511636 432612
rect 511670 432578 511726 432612
rect 511760 432578 511816 432612
rect 511850 432578 511906 432612
rect 511940 432578 511996 432612
rect 512030 432578 512082 432612
rect 511402 432522 512082 432578
rect 511402 432488 511456 432522
rect 511490 432488 511546 432522
rect 511580 432488 511636 432522
rect 511670 432488 511726 432522
rect 511760 432488 511816 432522
rect 511850 432488 511906 432522
rect 511940 432488 511996 432522
rect 512030 432488 512082 432522
rect 511402 432432 512082 432488
rect 511402 432398 511456 432432
rect 511490 432398 511546 432432
rect 511580 432398 511636 432432
rect 511670 432398 511726 432432
rect 511760 432398 511816 432432
rect 511850 432398 511906 432432
rect 511940 432398 511996 432432
rect 512030 432398 512082 432432
rect 511402 432346 512082 432398
rect 512690 432972 513370 433026
rect 512690 432938 512744 432972
rect 512778 432938 512834 432972
rect 512868 432938 512924 432972
rect 512958 432938 513014 432972
rect 513048 432938 513104 432972
rect 513138 432938 513194 432972
rect 513228 432938 513284 432972
rect 513318 432938 513370 432972
rect 512690 432882 513370 432938
rect 512690 432848 512744 432882
rect 512778 432848 512834 432882
rect 512868 432848 512924 432882
rect 512958 432848 513014 432882
rect 513048 432848 513104 432882
rect 513138 432848 513194 432882
rect 513228 432848 513284 432882
rect 513318 432848 513370 432882
rect 512690 432792 513370 432848
rect 512690 432758 512744 432792
rect 512778 432758 512834 432792
rect 512868 432758 512924 432792
rect 512958 432758 513014 432792
rect 513048 432758 513104 432792
rect 513138 432758 513194 432792
rect 513228 432758 513284 432792
rect 513318 432758 513370 432792
rect 512690 432702 513370 432758
rect 512690 432668 512744 432702
rect 512778 432668 512834 432702
rect 512868 432668 512924 432702
rect 512958 432668 513014 432702
rect 513048 432668 513104 432702
rect 513138 432668 513194 432702
rect 513228 432668 513284 432702
rect 513318 432668 513370 432702
rect 512690 432612 513370 432668
rect 512690 432578 512744 432612
rect 512778 432578 512834 432612
rect 512868 432578 512924 432612
rect 512958 432578 513014 432612
rect 513048 432578 513104 432612
rect 513138 432578 513194 432612
rect 513228 432578 513284 432612
rect 513318 432578 513370 432612
rect 512690 432522 513370 432578
rect 512690 432488 512744 432522
rect 512778 432488 512834 432522
rect 512868 432488 512924 432522
rect 512958 432488 513014 432522
rect 513048 432488 513104 432522
rect 513138 432488 513194 432522
rect 513228 432488 513284 432522
rect 513318 432488 513370 432522
rect 512690 432432 513370 432488
rect 512690 432398 512744 432432
rect 512778 432398 512834 432432
rect 512868 432398 512924 432432
rect 512958 432398 513014 432432
rect 513048 432398 513104 432432
rect 513138 432398 513194 432432
rect 513228 432398 513284 432432
rect 513318 432398 513370 432432
rect 512690 432346 513370 432398
rect 562258 455088 562316 455100
rect 562258 454112 562270 455088
rect 562304 454112 562316 455088
rect 562258 454100 562316 454112
rect 562516 455088 562574 455100
rect 562516 454112 562528 455088
rect 562562 454112 562574 455088
rect 562516 454100 562574 454112
rect 562774 455088 562832 455100
rect 562774 454112 562786 455088
rect 562820 454112 562832 455088
rect 562774 454100 562832 454112
rect 563032 455088 563090 455100
rect 563032 454112 563044 455088
rect 563078 454112 563090 455088
rect 563032 454100 563090 454112
rect 563290 455088 563348 455100
rect 563290 454112 563302 455088
rect 563336 454112 563348 455088
rect 563290 454100 563348 454112
rect 563548 455088 563606 455100
rect 563548 454112 563560 455088
rect 563594 454112 563606 455088
rect 563548 454100 563606 454112
rect 563806 455088 563864 455100
rect 563806 454112 563818 455088
rect 563852 454112 563864 455088
rect 563806 454100 563864 454112
rect 564064 455088 564122 455100
rect 564064 454112 564076 455088
rect 564110 454112 564122 455088
rect 564064 454100 564122 454112
rect 564322 455088 564380 455100
rect 564322 454112 564334 455088
rect 564368 454112 564380 455088
rect 564322 454100 564380 454112
rect 564580 455088 564638 455100
rect 564580 454112 564592 455088
rect 564626 454112 564638 455088
rect 564580 454100 564638 454112
rect 564838 455088 564896 455100
rect 564838 454112 564850 455088
rect 564884 454112 564896 455088
rect 564838 454100 564896 454112
rect 565096 455088 565154 455100
rect 565096 454112 565108 455088
rect 565142 454112 565154 455088
rect 565096 454100 565154 454112
rect 565354 455088 565412 455100
rect 565354 454112 565366 455088
rect 565400 454112 565412 455088
rect 565354 454100 565412 454112
rect 565612 455088 565670 455100
rect 565612 454112 565624 455088
rect 565658 454112 565670 455088
rect 565612 454100 565670 454112
rect 565870 455088 565928 455100
rect 565870 454112 565882 455088
rect 565916 454112 565928 455088
rect 565870 454100 565928 454112
rect 566128 455088 566186 455100
rect 566128 454112 566140 455088
rect 566174 454112 566186 455088
rect 566128 454100 566186 454112
rect 566386 455088 566444 455100
rect 566386 454112 566398 455088
rect 566432 454112 566444 455088
rect 566386 454100 566444 454112
rect 566644 455088 566702 455100
rect 566644 454112 566656 455088
rect 566690 454112 566702 455088
rect 566644 454100 566702 454112
rect 566902 455088 566960 455100
rect 566902 454112 566914 455088
rect 566948 454112 566960 455088
rect 566902 454100 566960 454112
rect 567160 455088 567218 455100
rect 567160 454112 567172 455088
rect 567206 454112 567218 455088
rect 567160 454100 567218 454112
rect 567418 455088 567476 455100
rect 567418 454112 567430 455088
rect 567464 454112 567476 455088
rect 567418 454100 567476 454112
<< ndiffc >>
rect 572430 494448 572464 495424
rect 572688 494448 572722 495424
rect 572946 494448 572980 495424
rect 573204 494448 573238 495424
rect 573462 494448 573496 495424
rect 573720 494448 573754 495424
rect 573978 494448 574012 495424
rect 574236 494448 574270 495424
rect 574494 494448 574528 495424
rect 574752 494448 574786 495424
rect 575010 494448 575044 495424
rect 575268 494448 575302 495424
rect 575526 494448 575560 495424
rect 575784 494448 575818 495424
rect 576042 494448 576076 495424
rect 576300 494448 576334 495424
rect 576558 494448 576592 495424
rect 576816 494448 576850 495424
rect 577074 494448 577108 495424
rect 577332 494448 577366 495424
rect 577590 494448 577624 495424
rect 506570 472730 506946 472764
rect 506570 472272 506946 472306
rect 506570 471814 506946 471848
rect 506570 471356 506946 471390
rect 506570 470898 506946 470932
rect 506570 470440 506946 470474
rect 506570 469982 506946 470016
rect 506292 467800 508068 467834
rect 506292 467342 508068 467376
rect 506292 467228 508068 467262
rect 506292 466770 508068 466804
rect 506292 466656 508068 466690
rect 506292 466198 508068 466232
rect 506292 466084 508068 466118
rect 506292 465626 508068 465660
rect 506292 465512 508068 465546
rect 506292 465054 508068 465088
rect 506292 464940 508068 464974
rect 506292 464482 508068 464516
rect 506292 464368 508068 464402
rect 506292 463910 508068 463944
rect 506292 463796 508068 463830
rect 506292 463338 508068 463372
rect 509786 462740 509820 468116
rect 510244 462740 510278 468116
rect 572430 454146 572464 455122
rect 572688 454146 572722 455122
rect 572946 454146 572980 455122
rect 573204 454146 573238 455122
rect 573462 454146 573496 455122
rect 573720 454146 573754 455122
rect 573978 454146 574012 455122
rect 574236 454146 574270 455122
rect 574494 454146 574528 455122
rect 574752 454146 574786 455122
rect 575010 454146 575044 455122
rect 575268 454146 575302 455122
rect 575526 454146 575560 455122
rect 575784 454146 575818 455122
rect 576042 454146 576076 455122
rect 576300 454146 576334 455122
rect 576558 454146 576592 455122
rect 576816 454146 576850 455122
rect 577074 454146 577108 455122
rect 577332 454146 577366 455122
rect 577590 454146 577624 455122
<< pdiffc >>
rect 562270 494414 562304 495390
rect 562528 494414 562562 495390
rect 562786 494414 562820 495390
rect 563044 494414 563078 495390
rect 563302 494414 563336 495390
rect 563560 494414 563594 495390
rect 563818 494414 563852 495390
rect 564076 494414 564110 495390
rect 564334 494414 564368 495390
rect 564592 494414 564626 495390
rect 564850 494414 564884 495390
rect 565108 494414 565142 495390
rect 565366 494414 565400 495390
rect 565624 494414 565658 495390
rect 565882 494414 565916 495390
rect 566140 494414 566174 495390
rect 566398 494414 566432 495390
rect 566656 494414 566690 495390
rect 566914 494414 566948 495390
rect 567172 494414 567206 495390
rect 567430 494414 567464 495390
rect 503100 469526 505656 469560
rect 503100 469068 505656 469102
rect 503100 468954 505656 468988
rect 503100 468496 505656 468530
rect 503100 468382 505656 468416
rect 503100 467924 505656 467958
rect 503100 467810 505656 467844
rect 503100 467352 505656 467386
rect 503100 467238 505656 467272
rect 503100 466780 505656 466814
rect 503100 466666 505656 466700
rect 503100 466208 505656 466242
rect 503100 466094 505656 466128
rect 503100 465636 505656 465670
rect 503100 465522 505656 465556
rect 503100 465064 505656 465098
rect 503100 464950 505656 464984
rect 503100 464492 505656 464526
rect 503100 464378 505656 464412
rect 503100 463920 505656 463954
rect 503100 463806 505656 463840
rect 503100 463348 505656 463382
rect 503100 463234 505656 463268
rect 503100 462776 505656 462810
rect 503100 462662 505656 462696
rect 503100 462204 505656 462238
rect 503100 462090 505656 462124
rect 503100 461632 505656 461666
rect 503138 459718 510854 459752
rect 503138 459260 510854 459294
rect 503138 458802 510854 458836
rect 503138 458344 510854 458378
rect 503138 457886 510854 457920
rect 503138 457428 510854 457462
rect 503138 456970 510854 457004
rect 503138 456512 510854 456546
rect 503138 456054 510854 456088
rect 503138 455596 510854 455630
rect 503138 455138 510854 455172
rect 503138 454680 510854 454714
rect 503138 453760 510854 453794
rect 503138 453302 510854 453336
rect 503138 452844 510854 452878
rect 503138 452386 510854 452420
rect 503138 451928 510854 451962
rect 503138 451470 510854 451504
rect 503138 451012 510854 451046
rect 503138 450554 510854 450588
rect 503138 450096 510854 450130
rect 503138 449638 510854 449672
rect 503138 449180 510854 449214
rect 503138 448260 510854 448294
rect 503138 447802 510854 447836
rect 503138 447344 510854 447378
rect 503138 446886 510854 446920
rect 503138 446428 510854 446462
rect 503138 445970 510854 446004
rect 503138 445512 510854 445546
rect 503138 445054 510854 445088
rect 503138 444596 510854 444630
rect 503138 444138 510854 444172
rect 503138 443680 510854 443714
rect 503138 443222 510854 443256
rect 503728 438090 503762 438124
rect 503818 438090 503852 438124
rect 503908 438090 503942 438124
rect 503998 438090 504032 438124
rect 504088 438090 504122 438124
rect 504178 438090 504212 438124
rect 504268 438090 504302 438124
rect 503728 438000 503762 438034
rect 503818 438000 503852 438034
rect 503908 438000 503942 438034
rect 503998 438000 504032 438034
rect 504088 438000 504122 438034
rect 504178 438000 504212 438034
rect 504268 438000 504302 438034
rect 503728 437910 503762 437944
rect 503818 437910 503852 437944
rect 503908 437910 503942 437944
rect 503998 437910 504032 437944
rect 504088 437910 504122 437944
rect 504178 437910 504212 437944
rect 504268 437910 504302 437944
rect 503728 437820 503762 437854
rect 503818 437820 503852 437854
rect 503908 437820 503942 437854
rect 503998 437820 504032 437854
rect 504088 437820 504122 437854
rect 504178 437820 504212 437854
rect 504268 437820 504302 437854
rect 503728 437730 503762 437764
rect 503818 437730 503852 437764
rect 503908 437730 503942 437764
rect 503998 437730 504032 437764
rect 504088 437730 504122 437764
rect 504178 437730 504212 437764
rect 504268 437730 504302 437764
rect 503728 437640 503762 437674
rect 503818 437640 503852 437674
rect 503908 437640 503942 437674
rect 503998 437640 504032 437674
rect 504088 437640 504122 437674
rect 504178 437640 504212 437674
rect 504268 437640 504302 437674
rect 503728 437550 503762 437584
rect 503818 437550 503852 437584
rect 503908 437550 503942 437584
rect 503998 437550 504032 437584
rect 504088 437550 504122 437584
rect 504178 437550 504212 437584
rect 504268 437550 504302 437584
rect 505016 438090 505050 438124
rect 505106 438090 505140 438124
rect 505196 438090 505230 438124
rect 505286 438090 505320 438124
rect 505376 438090 505410 438124
rect 505466 438090 505500 438124
rect 505556 438090 505590 438124
rect 505016 438000 505050 438034
rect 505106 438000 505140 438034
rect 505196 438000 505230 438034
rect 505286 438000 505320 438034
rect 505376 438000 505410 438034
rect 505466 438000 505500 438034
rect 505556 438000 505590 438034
rect 505016 437910 505050 437944
rect 505106 437910 505140 437944
rect 505196 437910 505230 437944
rect 505286 437910 505320 437944
rect 505376 437910 505410 437944
rect 505466 437910 505500 437944
rect 505556 437910 505590 437944
rect 505016 437820 505050 437854
rect 505106 437820 505140 437854
rect 505196 437820 505230 437854
rect 505286 437820 505320 437854
rect 505376 437820 505410 437854
rect 505466 437820 505500 437854
rect 505556 437820 505590 437854
rect 505016 437730 505050 437764
rect 505106 437730 505140 437764
rect 505196 437730 505230 437764
rect 505286 437730 505320 437764
rect 505376 437730 505410 437764
rect 505466 437730 505500 437764
rect 505556 437730 505590 437764
rect 505016 437640 505050 437674
rect 505106 437640 505140 437674
rect 505196 437640 505230 437674
rect 505286 437640 505320 437674
rect 505376 437640 505410 437674
rect 505466 437640 505500 437674
rect 505556 437640 505590 437674
rect 505016 437550 505050 437584
rect 505106 437550 505140 437584
rect 505196 437550 505230 437584
rect 505286 437550 505320 437584
rect 505376 437550 505410 437584
rect 505466 437550 505500 437584
rect 505556 437550 505590 437584
rect 506304 438090 506338 438124
rect 506394 438090 506428 438124
rect 506484 438090 506518 438124
rect 506574 438090 506608 438124
rect 506664 438090 506698 438124
rect 506754 438090 506788 438124
rect 506844 438090 506878 438124
rect 506304 438000 506338 438034
rect 506394 438000 506428 438034
rect 506484 438000 506518 438034
rect 506574 438000 506608 438034
rect 506664 438000 506698 438034
rect 506754 438000 506788 438034
rect 506844 438000 506878 438034
rect 506304 437910 506338 437944
rect 506394 437910 506428 437944
rect 506484 437910 506518 437944
rect 506574 437910 506608 437944
rect 506664 437910 506698 437944
rect 506754 437910 506788 437944
rect 506844 437910 506878 437944
rect 506304 437820 506338 437854
rect 506394 437820 506428 437854
rect 506484 437820 506518 437854
rect 506574 437820 506608 437854
rect 506664 437820 506698 437854
rect 506754 437820 506788 437854
rect 506844 437820 506878 437854
rect 506304 437730 506338 437764
rect 506394 437730 506428 437764
rect 506484 437730 506518 437764
rect 506574 437730 506608 437764
rect 506664 437730 506698 437764
rect 506754 437730 506788 437764
rect 506844 437730 506878 437764
rect 506304 437640 506338 437674
rect 506394 437640 506428 437674
rect 506484 437640 506518 437674
rect 506574 437640 506608 437674
rect 506664 437640 506698 437674
rect 506754 437640 506788 437674
rect 506844 437640 506878 437674
rect 506304 437550 506338 437584
rect 506394 437550 506428 437584
rect 506484 437550 506518 437584
rect 506574 437550 506608 437584
rect 506664 437550 506698 437584
rect 506754 437550 506788 437584
rect 506844 437550 506878 437584
rect 507592 438090 507626 438124
rect 507682 438090 507716 438124
rect 507772 438090 507806 438124
rect 507862 438090 507896 438124
rect 507952 438090 507986 438124
rect 508042 438090 508076 438124
rect 508132 438090 508166 438124
rect 507592 438000 507626 438034
rect 507682 438000 507716 438034
rect 507772 438000 507806 438034
rect 507862 438000 507896 438034
rect 507952 438000 507986 438034
rect 508042 438000 508076 438034
rect 508132 438000 508166 438034
rect 507592 437910 507626 437944
rect 507682 437910 507716 437944
rect 507772 437910 507806 437944
rect 507862 437910 507896 437944
rect 507952 437910 507986 437944
rect 508042 437910 508076 437944
rect 508132 437910 508166 437944
rect 507592 437820 507626 437854
rect 507682 437820 507716 437854
rect 507772 437820 507806 437854
rect 507862 437820 507896 437854
rect 507952 437820 507986 437854
rect 508042 437820 508076 437854
rect 508132 437820 508166 437854
rect 507592 437730 507626 437764
rect 507682 437730 507716 437764
rect 507772 437730 507806 437764
rect 507862 437730 507896 437764
rect 507952 437730 507986 437764
rect 508042 437730 508076 437764
rect 508132 437730 508166 437764
rect 507592 437640 507626 437674
rect 507682 437640 507716 437674
rect 507772 437640 507806 437674
rect 507862 437640 507896 437674
rect 507952 437640 507986 437674
rect 508042 437640 508076 437674
rect 508132 437640 508166 437674
rect 507592 437550 507626 437584
rect 507682 437550 507716 437584
rect 507772 437550 507806 437584
rect 507862 437550 507896 437584
rect 507952 437550 507986 437584
rect 508042 437550 508076 437584
rect 508132 437550 508166 437584
rect 508880 438090 508914 438124
rect 508970 438090 509004 438124
rect 509060 438090 509094 438124
rect 509150 438090 509184 438124
rect 509240 438090 509274 438124
rect 509330 438090 509364 438124
rect 509420 438090 509454 438124
rect 508880 438000 508914 438034
rect 508970 438000 509004 438034
rect 509060 438000 509094 438034
rect 509150 438000 509184 438034
rect 509240 438000 509274 438034
rect 509330 438000 509364 438034
rect 509420 438000 509454 438034
rect 508880 437910 508914 437944
rect 508970 437910 509004 437944
rect 509060 437910 509094 437944
rect 509150 437910 509184 437944
rect 509240 437910 509274 437944
rect 509330 437910 509364 437944
rect 509420 437910 509454 437944
rect 508880 437820 508914 437854
rect 508970 437820 509004 437854
rect 509060 437820 509094 437854
rect 509150 437820 509184 437854
rect 509240 437820 509274 437854
rect 509330 437820 509364 437854
rect 509420 437820 509454 437854
rect 508880 437730 508914 437764
rect 508970 437730 509004 437764
rect 509060 437730 509094 437764
rect 509150 437730 509184 437764
rect 509240 437730 509274 437764
rect 509330 437730 509364 437764
rect 509420 437730 509454 437764
rect 508880 437640 508914 437674
rect 508970 437640 509004 437674
rect 509060 437640 509094 437674
rect 509150 437640 509184 437674
rect 509240 437640 509274 437674
rect 509330 437640 509364 437674
rect 509420 437640 509454 437674
rect 508880 437550 508914 437584
rect 508970 437550 509004 437584
rect 509060 437550 509094 437584
rect 509150 437550 509184 437584
rect 509240 437550 509274 437584
rect 509330 437550 509364 437584
rect 509420 437550 509454 437584
rect 510168 438090 510202 438124
rect 510258 438090 510292 438124
rect 510348 438090 510382 438124
rect 510438 438090 510472 438124
rect 510528 438090 510562 438124
rect 510618 438090 510652 438124
rect 510708 438090 510742 438124
rect 510168 438000 510202 438034
rect 510258 438000 510292 438034
rect 510348 438000 510382 438034
rect 510438 438000 510472 438034
rect 510528 438000 510562 438034
rect 510618 438000 510652 438034
rect 510708 438000 510742 438034
rect 510168 437910 510202 437944
rect 510258 437910 510292 437944
rect 510348 437910 510382 437944
rect 510438 437910 510472 437944
rect 510528 437910 510562 437944
rect 510618 437910 510652 437944
rect 510708 437910 510742 437944
rect 510168 437820 510202 437854
rect 510258 437820 510292 437854
rect 510348 437820 510382 437854
rect 510438 437820 510472 437854
rect 510528 437820 510562 437854
rect 510618 437820 510652 437854
rect 510708 437820 510742 437854
rect 510168 437730 510202 437764
rect 510258 437730 510292 437764
rect 510348 437730 510382 437764
rect 510438 437730 510472 437764
rect 510528 437730 510562 437764
rect 510618 437730 510652 437764
rect 510708 437730 510742 437764
rect 510168 437640 510202 437674
rect 510258 437640 510292 437674
rect 510348 437640 510382 437674
rect 510438 437640 510472 437674
rect 510528 437640 510562 437674
rect 510618 437640 510652 437674
rect 510708 437640 510742 437674
rect 510168 437550 510202 437584
rect 510258 437550 510292 437584
rect 510348 437550 510382 437584
rect 510438 437550 510472 437584
rect 510528 437550 510562 437584
rect 510618 437550 510652 437584
rect 510708 437550 510742 437584
rect 511456 438090 511490 438124
rect 511546 438090 511580 438124
rect 511636 438090 511670 438124
rect 511726 438090 511760 438124
rect 511816 438090 511850 438124
rect 511906 438090 511940 438124
rect 511996 438090 512030 438124
rect 511456 438000 511490 438034
rect 511546 438000 511580 438034
rect 511636 438000 511670 438034
rect 511726 438000 511760 438034
rect 511816 438000 511850 438034
rect 511906 438000 511940 438034
rect 511996 438000 512030 438034
rect 511456 437910 511490 437944
rect 511546 437910 511580 437944
rect 511636 437910 511670 437944
rect 511726 437910 511760 437944
rect 511816 437910 511850 437944
rect 511906 437910 511940 437944
rect 511996 437910 512030 437944
rect 511456 437820 511490 437854
rect 511546 437820 511580 437854
rect 511636 437820 511670 437854
rect 511726 437820 511760 437854
rect 511816 437820 511850 437854
rect 511906 437820 511940 437854
rect 511996 437820 512030 437854
rect 511456 437730 511490 437764
rect 511546 437730 511580 437764
rect 511636 437730 511670 437764
rect 511726 437730 511760 437764
rect 511816 437730 511850 437764
rect 511906 437730 511940 437764
rect 511996 437730 512030 437764
rect 511456 437640 511490 437674
rect 511546 437640 511580 437674
rect 511636 437640 511670 437674
rect 511726 437640 511760 437674
rect 511816 437640 511850 437674
rect 511906 437640 511940 437674
rect 511996 437640 512030 437674
rect 511456 437550 511490 437584
rect 511546 437550 511580 437584
rect 511636 437550 511670 437584
rect 511726 437550 511760 437584
rect 511816 437550 511850 437584
rect 511906 437550 511940 437584
rect 511996 437550 512030 437584
rect 512744 438090 512778 438124
rect 512834 438090 512868 438124
rect 512924 438090 512958 438124
rect 513014 438090 513048 438124
rect 513104 438090 513138 438124
rect 513194 438090 513228 438124
rect 513284 438090 513318 438124
rect 512744 438000 512778 438034
rect 512834 438000 512868 438034
rect 512924 438000 512958 438034
rect 513014 438000 513048 438034
rect 513104 438000 513138 438034
rect 513194 438000 513228 438034
rect 513284 438000 513318 438034
rect 512744 437910 512778 437944
rect 512834 437910 512868 437944
rect 512924 437910 512958 437944
rect 513014 437910 513048 437944
rect 513104 437910 513138 437944
rect 513194 437910 513228 437944
rect 513284 437910 513318 437944
rect 512744 437820 512778 437854
rect 512834 437820 512868 437854
rect 512924 437820 512958 437854
rect 513014 437820 513048 437854
rect 513104 437820 513138 437854
rect 513194 437820 513228 437854
rect 513284 437820 513318 437854
rect 512744 437730 512778 437764
rect 512834 437730 512868 437764
rect 512924 437730 512958 437764
rect 513014 437730 513048 437764
rect 513104 437730 513138 437764
rect 513194 437730 513228 437764
rect 513284 437730 513318 437764
rect 512744 437640 512778 437674
rect 512834 437640 512868 437674
rect 512924 437640 512958 437674
rect 513014 437640 513048 437674
rect 513104 437640 513138 437674
rect 513194 437640 513228 437674
rect 513284 437640 513318 437674
rect 512744 437550 512778 437584
rect 512834 437550 512868 437584
rect 512924 437550 512958 437584
rect 513014 437550 513048 437584
rect 513104 437550 513138 437584
rect 513194 437550 513228 437584
rect 513284 437550 513318 437584
rect 503728 436802 503762 436836
rect 503818 436802 503852 436836
rect 503908 436802 503942 436836
rect 503998 436802 504032 436836
rect 504088 436802 504122 436836
rect 504178 436802 504212 436836
rect 504268 436802 504302 436836
rect 503728 436712 503762 436746
rect 503818 436712 503852 436746
rect 503908 436712 503942 436746
rect 503998 436712 504032 436746
rect 504088 436712 504122 436746
rect 504178 436712 504212 436746
rect 504268 436712 504302 436746
rect 503728 436622 503762 436656
rect 503818 436622 503852 436656
rect 503908 436622 503942 436656
rect 503998 436622 504032 436656
rect 504088 436622 504122 436656
rect 504178 436622 504212 436656
rect 504268 436622 504302 436656
rect 503728 436532 503762 436566
rect 503818 436532 503852 436566
rect 503908 436532 503942 436566
rect 503998 436532 504032 436566
rect 504088 436532 504122 436566
rect 504178 436532 504212 436566
rect 504268 436532 504302 436566
rect 503728 436442 503762 436476
rect 503818 436442 503852 436476
rect 503908 436442 503942 436476
rect 503998 436442 504032 436476
rect 504088 436442 504122 436476
rect 504178 436442 504212 436476
rect 504268 436442 504302 436476
rect 503728 436352 503762 436386
rect 503818 436352 503852 436386
rect 503908 436352 503942 436386
rect 503998 436352 504032 436386
rect 504088 436352 504122 436386
rect 504178 436352 504212 436386
rect 504268 436352 504302 436386
rect 503728 436262 503762 436296
rect 503818 436262 503852 436296
rect 503908 436262 503942 436296
rect 503998 436262 504032 436296
rect 504088 436262 504122 436296
rect 504178 436262 504212 436296
rect 504268 436262 504302 436296
rect 505016 436802 505050 436836
rect 505106 436802 505140 436836
rect 505196 436802 505230 436836
rect 505286 436802 505320 436836
rect 505376 436802 505410 436836
rect 505466 436802 505500 436836
rect 505556 436802 505590 436836
rect 505016 436712 505050 436746
rect 505106 436712 505140 436746
rect 505196 436712 505230 436746
rect 505286 436712 505320 436746
rect 505376 436712 505410 436746
rect 505466 436712 505500 436746
rect 505556 436712 505590 436746
rect 505016 436622 505050 436656
rect 505106 436622 505140 436656
rect 505196 436622 505230 436656
rect 505286 436622 505320 436656
rect 505376 436622 505410 436656
rect 505466 436622 505500 436656
rect 505556 436622 505590 436656
rect 505016 436532 505050 436566
rect 505106 436532 505140 436566
rect 505196 436532 505230 436566
rect 505286 436532 505320 436566
rect 505376 436532 505410 436566
rect 505466 436532 505500 436566
rect 505556 436532 505590 436566
rect 505016 436442 505050 436476
rect 505106 436442 505140 436476
rect 505196 436442 505230 436476
rect 505286 436442 505320 436476
rect 505376 436442 505410 436476
rect 505466 436442 505500 436476
rect 505556 436442 505590 436476
rect 505016 436352 505050 436386
rect 505106 436352 505140 436386
rect 505196 436352 505230 436386
rect 505286 436352 505320 436386
rect 505376 436352 505410 436386
rect 505466 436352 505500 436386
rect 505556 436352 505590 436386
rect 505016 436262 505050 436296
rect 505106 436262 505140 436296
rect 505196 436262 505230 436296
rect 505286 436262 505320 436296
rect 505376 436262 505410 436296
rect 505466 436262 505500 436296
rect 505556 436262 505590 436296
rect 506304 436802 506338 436836
rect 506394 436802 506428 436836
rect 506484 436802 506518 436836
rect 506574 436802 506608 436836
rect 506664 436802 506698 436836
rect 506754 436802 506788 436836
rect 506844 436802 506878 436836
rect 506304 436712 506338 436746
rect 506394 436712 506428 436746
rect 506484 436712 506518 436746
rect 506574 436712 506608 436746
rect 506664 436712 506698 436746
rect 506754 436712 506788 436746
rect 506844 436712 506878 436746
rect 506304 436622 506338 436656
rect 506394 436622 506428 436656
rect 506484 436622 506518 436656
rect 506574 436622 506608 436656
rect 506664 436622 506698 436656
rect 506754 436622 506788 436656
rect 506844 436622 506878 436656
rect 506304 436532 506338 436566
rect 506394 436532 506428 436566
rect 506484 436532 506518 436566
rect 506574 436532 506608 436566
rect 506664 436532 506698 436566
rect 506754 436532 506788 436566
rect 506844 436532 506878 436566
rect 506304 436442 506338 436476
rect 506394 436442 506428 436476
rect 506484 436442 506518 436476
rect 506574 436442 506608 436476
rect 506664 436442 506698 436476
rect 506754 436442 506788 436476
rect 506844 436442 506878 436476
rect 506304 436352 506338 436386
rect 506394 436352 506428 436386
rect 506484 436352 506518 436386
rect 506574 436352 506608 436386
rect 506664 436352 506698 436386
rect 506754 436352 506788 436386
rect 506844 436352 506878 436386
rect 506304 436262 506338 436296
rect 506394 436262 506428 436296
rect 506484 436262 506518 436296
rect 506574 436262 506608 436296
rect 506664 436262 506698 436296
rect 506754 436262 506788 436296
rect 506844 436262 506878 436296
rect 507592 436802 507626 436836
rect 507682 436802 507716 436836
rect 507772 436802 507806 436836
rect 507862 436802 507896 436836
rect 507952 436802 507986 436836
rect 508042 436802 508076 436836
rect 508132 436802 508166 436836
rect 507592 436712 507626 436746
rect 507682 436712 507716 436746
rect 507772 436712 507806 436746
rect 507862 436712 507896 436746
rect 507952 436712 507986 436746
rect 508042 436712 508076 436746
rect 508132 436712 508166 436746
rect 507592 436622 507626 436656
rect 507682 436622 507716 436656
rect 507772 436622 507806 436656
rect 507862 436622 507896 436656
rect 507952 436622 507986 436656
rect 508042 436622 508076 436656
rect 508132 436622 508166 436656
rect 507592 436532 507626 436566
rect 507682 436532 507716 436566
rect 507772 436532 507806 436566
rect 507862 436532 507896 436566
rect 507952 436532 507986 436566
rect 508042 436532 508076 436566
rect 508132 436532 508166 436566
rect 507592 436442 507626 436476
rect 507682 436442 507716 436476
rect 507772 436442 507806 436476
rect 507862 436442 507896 436476
rect 507952 436442 507986 436476
rect 508042 436442 508076 436476
rect 508132 436442 508166 436476
rect 507592 436352 507626 436386
rect 507682 436352 507716 436386
rect 507772 436352 507806 436386
rect 507862 436352 507896 436386
rect 507952 436352 507986 436386
rect 508042 436352 508076 436386
rect 508132 436352 508166 436386
rect 507592 436262 507626 436296
rect 507682 436262 507716 436296
rect 507772 436262 507806 436296
rect 507862 436262 507896 436296
rect 507952 436262 507986 436296
rect 508042 436262 508076 436296
rect 508132 436262 508166 436296
rect 508880 436802 508914 436836
rect 508970 436802 509004 436836
rect 509060 436802 509094 436836
rect 509150 436802 509184 436836
rect 509240 436802 509274 436836
rect 509330 436802 509364 436836
rect 509420 436802 509454 436836
rect 508880 436712 508914 436746
rect 508970 436712 509004 436746
rect 509060 436712 509094 436746
rect 509150 436712 509184 436746
rect 509240 436712 509274 436746
rect 509330 436712 509364 436746
rect 509420 436712 509454 436746
rect 508880 436622 508914 436656
rect 508970 436622 509004 436656
rect 509060 436622 509094 436656
rect 509150 436622 509184 436656
rect 509240 436622 509274 436656
rect 509330 436622 509364 436656
rect 509420 436622 509454 436656
rect 508880 436532 508914 436566
rect 508970 436532 509004 436566
rect 509060 436532 509094 436566
rect 509150 436532 509184 436566
rect 509240 436532 509274 436566
rect 509330 436532 509364 436566
rect 509420 436532 509454 436566
rect 508880 436442 508914 436476
rect 508970 436442 509004 436476
rect 509060 436442 509094 436476
rect 509150 436442 509184 436476
rect 509240 436442 509274 436476
rect 509330 436442 509364 436476
rect 509420 436442 509454 436476
rect 508880 436352 508914 436386
rect 508970 436352 509004 436386
rect 509060 436352 509094 436386
rect 509150 436352 509184 436386
rect 509240 436352 509274 436386
rect 509330 436352 509364 436386
rect 509420 436352 509454 436386
rect 508880 436262 508914 436296
rect 508970 436262 509004 436296
rect 509060 436262 509094 436296
rect 509150 436262 509184 436296
rect 509240 436262 509274 436296
rect 509330 436262 509364 436296
rect 509420 436262 509454 436296
rect 510168 436802 510202 436836
rect 510258 436802 510292 436836
rect 510348 436802 510382 436836
rect 510438 436802 510472 436836
rect 510528 436802 510562 436836
rect 510618 436802 510652 436836
rect 510708 436802 510742 436836
rect 510168 436712 510202 436746
rect 510258 436712 510292 436746
rect 510348 436712 510382 436746
rect 510438 436712 510472 436746
rect 510528 436712 510562 436746
rect 510618 436712 510652 436746
rect 510708 436712 510742 436746
rect 510168 436622 510202 436656
rect 510258 436622 510292 436656
rect 510348 436622 510382 436656
rect 510438 436622 510472 436656
rect 510528 436622 510562 436656
rect 510618 436622 510652 436656
rect 510708 436622 510742 436656
rect 510168 436532 510202 436566
rect 510258 436532 510292 436566
rect 510348 436532 510382 436566
rect 510438 436532 510472 436566
rect 510528 436532 510562 436566
rect 510618 436532 510652 436566
rect 510708 436532 510742 436566
rect 510168 436442 510202 436476
rect 510258 436442 510292 436476
rect 510348 436442 510382 436476
rect 510438 436442 510472 436476
rect 510528 436442 510562 436476
rect 510618 436442 510652 436476
rect 510708 436442 510742 436476
rect 510168 436352 510202 436386
rect 510258 436352 510292 436386
rect 510348 436352 510382 436386
rect 510438 436352 510472 436386
rect 510528 436352 510562 436386
rect 510618 436352 510652 436386
rect 510708 436352 510742 436386
rect 510168 436262 510202 436296
rect 510258 436262 510292 436296
rect 510348 436262 510382 436296
rect 510438 436262 510472 436296
rect 510528 436262 510562 436296
rect 510618 436262 510652 436296
rect 510708 436262 510742 436296
rect 511456 436802 511490 436836
rect 511546 436802 511580 436836
rect 511636 436802 511670 436836
rect 511726 436802 511760 436836
rect 511816 436802 511850 436836
rect 511906 436802 511940 436836
rect 511996 436802 512030 436836
rect 511456 436712 511490 436746
rect 511546 436712 511580 436746
rect 511636 436712 511670 436746
rect 511726 436712 511760 436746
rect 511816 436712 511850 436746
rect 511906 436712 511940 436746
rect 511996 436712 512030 436746
rect 511456 436622 511490 436656
rect 511546 436622 511580 436656
rect 511636 436622 511670 436656
rect 511726 436622 511760 436656
rect 511816 436622 511850 436656
rect 511906 436622 511940 436656
rect 511996 436622 512030 436656
rect 511456 436532 511490 436566
rect 511546 436532 511580 436566
rect 511636 436532 511670 436566
rect 511726 436532 511760 436566
rect 511816 436532 511850 436566
rect 511906 436532 511940 436566
rect 511996 436532 512030 436566
rect 511456 436442 511490 436476
rect 511546 436442 511580 436476
rect 511636 436442 511670 436476
rect 511726 436442 511760 436476
rect 511816 436442 511850 436476
rect 511906 436442 511940 436476
rect 511996 436442 512030 436476
rect 511456 436352 511490 436386
rect 511546 436352 511580 436386
rect 511636 436352 511670 436386
rect 511726 436352 511760 436386
rect 511816 436352 511850 436386
rect 511906 436352 511940 436386
rect 511996 436352 512030 436386
rect 511456 436262 511490 436296
rect 511546 436262 511580 436296
rect 511636 436262 511670 436296
rect 511726 436262 511760 436296
rect 511816 436262 511850 436296
rect 511906 436262 511940 436296
rect 511996 436262 512030 436296
rect 512744 436802 512778 436836
rect 512834 436802 512868 436836
rect 512924 436802 512958 436836
rect 513014 436802 513048 436836
rect 513104 436802 513138 436836
rect 513194 436802 513228 436836
rect 513284 436802 513318 436836
rect 512744 436712 512778 436746
rect 512834 436712 512868 436746
rect 512924 436712 512958 436746
rect 513014 436712 513048 436746
rect 513104 436712 513138 436746
rect 513194 436712 513228 436746
rect 513284 436712 513318 436746
rect 512744 436622 512778 436656
rect 512834 436622 512868 436656
rect 512924 436622 512958 436656
rect 513014 436622 513048 436656
rect 513104 436622 513138 436656
rect 513194 436622 513228 436656
rect 513284 436622 513318 436656
rect 512744 436532 512778 436566
rect 512834 436532 512868 436566
rect 512924 436532 512958 436566
rect 513014 436532 513048 436566
rect 513104 436532 513138 436566
rect 513194 436532 513228 436566
rect 513284 436532 513318 436566
rect 512744 436442 512778 436476
rect 512834 436442 512868 436476
rect 512924 436442 512958 436476
rect 513014 436442 513048 436476
rect 513104 436442 513138 436476
rect 513194 436442 513228 436476
rect 513284 436442 513318 436476
rect 512744 436352 512778 436386
rect 512834 436352 512868 436386
rect 512924 436352 512958 436386
rect 513014 436352 513048 436386
rect 513104 436352 513138 436386
rect 513194 436352 513228 436386
rect 513284 436352 513318 436386
rect 512744 436262 512778 436296
rect 512834 436262 512868 436296
rect 512924 436262 512958 436296
rect 513014 436262 513048 436296
rect 513104 436262 513138 436296
rect 513194 436262 513228 436296
rect 513284 436262 513318 436296
rect 503728 435514 503762 435548
rect 503818 435514 503852 435548
rect 503908 435514 503942 435548
rect 503998 435514 504032 435548
rect 504088 435514 504122 435548
rect 504178 435514 504212 435548
rect 504268 435514 504302 435548
rect 503728 435424 503762 435458
rect 503818 435424 503852 435458
rect 503908 435424 503942 435458
rect 503998 435424 504032 435458
rect 504088 435424 504122 435458
rect 504178 435424 504212 435458
rect 504268 435424 504302 435458
rect 503728 435334 503762 435368
rect 503818 435334 503852 435368
rect 503908 435334 503942 435368
rect 503998 435334 504032 435368
rect 504088 435334 504122 435368
rect 504178 435334 504212 435368
rect 504268 435334 504302 435368
rect 503728 435244 503762 435278
rect 503818 435244 503852 435278
rect 503908 435244 503942 435278
rect 503998 435244 504032 435278
rect 504088 435244 504122 435278
rect 504178 435244 504212 435278
rect 504268 435244 504302 435278
rect 503728 435154 503762 435188
rect 503818 435154 503852 435188
rect 503908 435154 503942 435188
rect 503998 435154 504032 435188
rect 504088 435154 504122 435188
rect 504178 435154 504212 435188
rect 504268 435154 504302 435188
rect 503728 435064 503762 435098
rect 503818 435064 503852 435098
rect 503908 435064 503942 435098
rect 503998 435064 504032 435098
rect 504088 435064 504122 435098
rect 504178 435064 504212 435098
rect 504268 435064 504302 435098
rect 503728 434974 503762 435008
rect 503818 434974 503852 435008
rect 503908 434974 503942 435008
rect 503998 434974 504032 435008
rect 504088 434974 504122 435008
rect 504178 434974 504212 435008
rect 504268 434974 504302 435008
rect 505016 435514 505050 435548
rect 505106 435514 505140 435548
rect 505196 435514 505230 435548
rect 505286 435514 505320 435548
rect 505376 435514 505410 435548
rect 505466 435514 505500 435548
rect 505556 435514 505590 435548
rect 505016 435424 505050 435458
rect 505106 435424 505140 435458
rect 505196 435424 505230 435458
rect 505286 435424 505320 435458
rect 505376 435424 505410 435458
rect 505466 435424 505500 435458
rect 505556 435424 505590 435458
rect 505016 435334 505050 435368
rect 505106 435334 505140 435368
rect 505196 435334 505230 435368
rect 505286 435334 505320 435368
rect 505376 435334 505410 435368
rect 505466 435334 505500 435368
rect 505556 435334 505590 435368
rect 505016 435244 505050 435278
rect 505106 435244 505140 435278
rect 505196 435244 505230 435278
rect 505286 435244 505320 435278
rect 505376 435244 505410 435278
rect 505466 435244 505500 435278
rect 505556 435244 505590 435278
rect 505016 435154 505050 435188
rect 505106 435154 505140 435188
rect 505196 435154 505230 435188
rect 505286 435154 505320 435188
rect 505376 435154 505410 435188
rect 505466 435154 505500 435188
rect 505556 435154 505590 435188
rect 505016 435064 505050 435098
rect 505106 435064 505140 435098
rect 505196 435064 505230 435098
rect 505286 435064 505320 435098
rect 505376 435064 505410 435098
rect 505466 435064 505500 435098
rect 505556 435064 505590 435098
rect 505016 434974 505050 435008
rect 505106 434974 505140 435008
rect 505196 434974 505230 435008
rect 505286 434974 505320 435008
rect 505376 434974 505410 435008
rect 505466 434974 505500 435008
rect 505556 434974 505590 435008
rect 506304 435514 506338 435548
rect 506394 435514 506428 435548
rect 506484 435514 506518 435548
rect 506574 435514 506608 435548
rect 506664 435514 506698 435548
rect 506754 435514 506788 435548
rect 506844 435514 506878 435548
rect 506304 435424 506338 435458
rect 506394 435424 506428 435458
rect 506484 435424 506518 435458
rect 506574 435424 506608 435458
rect 506664 435424 506698 435458
rect 506754 435424 506788 435458
rect 506844 435424 506878 435458
rect 506304 435334 506338 435368
rect 506394 435334 506428 435368
rect 506484 435334 506518 435368
rect 506574 435334 506608 435368
rect 506664 435334 506698 435368
rect 506754 435334 506788 435368
rect 506844 435334 506878 435368
rect 506304 435244 506338 435278
rect 506394 435244 506428 435278
rect 506484 435244 506518 435278
rect 506574 435244 506608 435278
rect 506664 435244 506698 435278
rect 506754 435244 506788 435278
rect 506844 435244 506878 435278
rect 506304 435154 506338 435188
rect 506394 435154 506428 435188
rect 506484 435154 506518 435188
rect 506574 435154 506608 435188
rect 506664 435154 506698 435188
rect 506754 435154 506788 435188
rect 506844 435154 506878 435188
rect 506304 435064 506338 435098
rect 506394 435064 506428 435098
rect 506484 435064 506518 435098
rect 506574 435064 506608 435098
rect 506664 435064 506698 435098
rect 506754 435064 506788 435098
rect 506844 435064 506878 435098
rect 506304 434974 506338 435008
rect 506394 434974 506428 435008
rect 506484 434974 506518 435008
rect 506574 434974 506608 435008
rect 506664 434974 506698 435008
rect 506754 434974 506788 435008
rect 506844 434974 506878 435008
rect 507592 435514 507626 435548
rect 507682 435514 507716 435548
rect 507772 435514 507806 435548
rect 507862 435514 507896 435548
rect 507952 435514 507986 435548
rect 508042 435514 508076 435548
rect 508132 435514 508166 435548
rect 507592 435424 507626 435458
rect 507682 435424 507716 435458
rect 507772 435424 507806 435458
rect 507862 435424 507896 435458
rect 507952 435424 507986 435458
rect 508042 435424 508076 435458
rect 508132 435424 508166 435458
rect 507592 435334 507626 435368
rect 507682 435334 507716 435368
rect 507772 435334 507806 435368
rect 507862 435334 507896 435368
rect 507952 435334 507986 435368
rect 508042 435334 508076 435368
rect 508132 435334 508166 435368
rect 507592 435244 507626 435278
rect 507682 435244 507716 435278
rect 507772 435244 507806 435278
rect 507862 435244 507896 435278
rect 507952 435244 507986 435278
rect 508042 435244 508076 435278
rect 508132 435244 508166 435278
rect 507592 435154 507626 435188
rect 507682 435154 507716 435188
rect 507772 435154 507806 435188
rect 507862 435154 507896 435188
rect 507952 435154 507986 435188
rect 508042 435154 508076 435188
rect 508132 435154 508166 435188
rect 507592 435064 507626 435098
rect 507682 435064 507716 435098
rect 507772 435064 507806 435098
rect 507862 435064 507896 435098
rect 507952 435064 507986 435098
rect 508042 435064 508076 435098
rect 508132 435064 508166 435098
rect 507592 434974 507626 435008
rect 507682 434974 507716 435008
rect 507772 434974 507806 435008
rect 507862 434974 507896 435008
rect 507952 434974 507986 435008
rect 508042 434974 508076 435008
rect 508132 434974 508166 435008
rect 508880 435514 508914 435548
rect 508970 435514 509004 435548
rect 509060 435514 509094 435548
rect 509150 435514 509184 435548
rect 509240 435514 509274 435548
rect 509330 435514 509364 435548
rect 509420 435514 509454 435548
rect 508880 435424 508914 435458
rect 508970 435424 509004 435458
rect 509060 435424 509094 435458
rect 509150 435424 509184 435458
rect 509240 435424 509274 435458
rect 509330 435424 509364 435458
rect 509420 435424 509454 435458
rect 508880 435334 508914 435368
rect 508970 435334 509004 435368
rect 509060 435334 509094 435368
rect 509150 435334 509184 435368
rect 509240 435334 509274 435368
rect 509330 435334 509364 435368
rect 509420 435334 509454 435368
rect 508880 435244 508914 435278
rect 508970 435244 509004 435278
rect 509060 435244 509094 435278
rect 509150 435244 509184 435278
rect 509240 435244 509274 435278
rect 509330 435244 509364 435278
rect 509420 435244 509454 435278
rect 508880 435154 508914 435188
rect 508970 435154 509004 435188
rect 509060 435154 509094 435188
rect 509150 435154 509184 435188
rect 509240 435154 509274 435188
rect 509330 435154 509364 435188
rect 509420 435154 509454 435188
rect 508880 435064 508914 435098
rect 508970 435064 509004 435098
rect 509060 435064 509094 435098
rect 509150 435064 509184 435098
rect 509240 435064 509274 435098
rect 509330 435064 509364 435098
rect 509420 435064 509454 435098
rect 508880 434974 508914 435008
rect 508970 434974 509004 435008
rect 509060 434974 509094 435008
rect 509150 434974 509184 435008
rect 509240 434974 509274 435008
rect 509330 434974 509364 435008
rect 509420 434974 509454 435008
rect 510168 435514 510202 435548
rect 510258 435514 510292 435548
rect 510348 435514 510382 435548
rect 510438 435514 510472 435548
rect 510528 435514 510562 435548
rect 510618 435514 510652 435548
rect 510708 435514 510742 435548
rect 510168 435424 510202 435458
rect 510258 435424 510292 435458
rect 510348 435424 510382 435458
rect 510438 435424 510472 435458
rect 510528 435424 510562 435458
rect 510618 435424 510652 435458
rect 510708 435424 510742 435458
rect 510168 435334 510202 435368
rect 510258 435334 510292 435368
rect 510348 435334 510382 435368
rect 510438 435334 510472 435368
rect 510528 435334 510562 435368
rect 510618 435334 510652 435368
rect 510708 435334 510742 435368
rect 510168 435244 510202 435278
rect 510258 435244 510292 435278
rect 510348 435244 510382 435278
rect 510438 435244 510472 435278
rect 510528 435244 510562 435278
rect 510618 435244 510652 435278
rect 510708 435244 510742 435278
rect 510168 435154 510202 435188
rect 510258 435154 510292 435188
rect 510348 435154 510382 435188
rect 510438 435154 510472 435188
rect 510528 435154 510562 435188
rect 510618 435154 510652 435188
rect 510708 435154 510742 435188
rect 510168 435064 510202 435098
rect 510258 435064 510292 435098
rect 510348 435064 510382 435098
rect 510438 435064 510472 435098
rect 510528 435064 510562 435098
rect 510618 435064 510652 435098
rect 510708 435064 510742 435098
rect 510168 434974 510202 435008
rect 510258 434974 510292 435008
rect 510348 434974 510382 435008
rect 510438 434974 510472 435008
rect 510528 434974 510562 435008
rect 510618 434974 510652 435008
rect 510708 434974 510742 435008
rect 511456 435514 511490 435548
rect 511546 435514 511580 435548
rect 511636 435514 511670 435548
rect 511726 435514 511760 435548
rect 511816 435514 511850 435548
rect 511906 435514 511940 435548
rect 511996 435514 512030 435548
rect 511456 435424 511490 435458
rect 511546 435424 511580 435458
rect 511636 435424 511670 435458
rect 511726 435424 511760 435458
rect 511816 435424 511850 435458
rect 511906 435424 511940 435458
rect 511996 435424 512030 435458
rect 511456 435334 511490 435368
rect 511546 435334 511580 435368
rect 511636 435334 511670 435368
rect 511726 435334 511760 435368
rect 511816 435334 511850 435368
rect 511906 435334 511940 435368
rect 511996 435334 512030 435368
rect 511456 435244 511490 435278
rect 511546 435244 511580 435278
rect 511636 435244 511670 435278
rect 511726 435244 511760 435278
rect 511816 435244 511850 435278
rect 511906 435244 511940 435278
rect 511996 435244 512030 435278
rect 511456 435154 511490 435188
rect 511546 435154 511580 435188
rect 511636 435154 511670 435188
rect 511726 435154 511760 435188
rect 511816 435154 511850 435188
rect 511906 435154 511940 435188
rect 511996 435154 512030 435188
rect 511456 435064 511490 435098
rect 511546 435064 511580 435098
rect 511636 435064 511670 435098
rect 511726 435064 511760 435098
rect 511816 435064 511850 435098
rect 511906 435064 511940 435098
rect 511996 435064 512030 435098
rect 511456 434974 511490 435008
rect 511546 434974 511580 435008
rect 511636 434974 511670 435008
rect 511726 434974 511760 435008
rect 511816 434974 511850 435008
rect 511906 434974 511940 435008
rect 511996 434974 512030 435008
rect 512744 435514 512778 435548
rect 512834 435514 512868 435548
rect 512924 435514 512958 435548
rect 513014 435514 513048 435548
rect 513104 435514 513138 435548
rect 513194 435514 513228 435548
rect 513284 435514 513318 435548
rect 512744 435424 512778 435458
rect 512834 435424 512868 435458
rect 512924 435424 512958 435458
rect 513014 435424 513048 435458
rect 513104 435424 513138 435458
rect 513194 435424 513228 435458
rect 513284 435424 513318 435458
rect 512744 435334 512778 435368
rect 512834 435334 512868 435368
rect 512924 435334 512958 435368
rect 513014 435334 513048 435368
rect 513104 435334 513138 435368
rect 513194 435334 513228 435368
rect 513284 435334 513318 435368
rect 512744 435244 512778 435278
rect 512834 435244 512868 435278
rect 512924 435244 512958 435278
rect 513014 435244 513048 435278
rect 513104 435244 513138 435278
rect 513194 435244 513228 435278
rect 513284 435244 513318 435278
rect 512744 435154 512778 435188
rect 512834 435154 512868 435188
rect 512924 435154 512958 435188
rect 513014 435154 513048 435188
rect 513104 435154 513138 435188
rect 513194 435154 513228 435188
rect 513284 435154 513318 435188
rect 512744 435064 512778 435098
rect 512834 435064 512868 435098
rect 512924 435064 512958 435098
rect 513014 435064 513048 435098
rect 513104 435064 513138 435098
rect 513194 435064 513228 435098
rect 513284 435064 513318 435098
rect 512744 434974 512778 435008
rect 512834 434974 512868 435008
rect 512924 434974 512958 435008
rect 513014 434974 513048 435008
rect 513104 434974 513138 435008
rect 513194 434974 513228 435008
rect 513284 434974 513318 435008
rect 503728 434226 503762 434260
rect 503818 434226 503852 434260
rect 503908 434226 503942 434260
rect 503998 434226 504032 434260
rect 504088 434226 504122 434260
rect 504178 434226 504212 434260
rect 504268 434226 504302 434260
rect 503728 434136 503762 434170
rect 503818 434136 503852 434170
rect 503908 434136 503942 434170
rect 503998 434136 504032 434170
rect 504088 434136 504122 434170
rect 504178 434136 504212 434170
rect 504268 434136 504302 434170
rect 503728 434046 503762 434080
rect 503818 434046 503852 434080
rect 503908 434046 503942 434080
rect 503998 434046 504032 434080
rect 504088 434046 504122 434080
rect 504178 434046 504212 434080
rect 504268 434046 504302 434080
rect 503728 433956 503762 433990
rect 503818 433956 503852 433990
rect 503908 433956 503942 433990
rect 503998 433956 504032 433990
rect 504088 433956 504122 433990
rect 504178 433956 504212 433990
rect 504268 433956 504302 433990
rect 503728 433866 503762 433900
rect 503818 433866 503852 433900
rect 503908 433866 503942 433900
rect 503998 433866 504032 433900
rect 504088 433866 504122 433900
rect 504178 433866 504212 433900
rect 504268 433866 504302 433900
rect 503728 433776 503762 433810
rect 503818 433776 503852 433810
rect 503908 433776 503942 433810
rect 503998 433776 504032 433810
rect 504088 433776 504122 433810
rect 504178 433776 504212 433810
rect 504268 433776 504302 433810
rect 503728 433686 503762 433720
rect 503818 433686 503852 433720
rect 503908 433686 503942 433720
rect 503998 433686 504032 433720
rect 504088 433686 504122 433720
rect 504178 433686 504212 433720
rect 504268 433686 504302 433720
rect 505016 434226 505050 434260
rect 505106 434226 505140 434260
rect 505196 434226 505230 434260
rect 505286 434226 505320 434260
rect 505376 434226 505410 434260
rect 505466 434226 505500 434260
rect 505556 434226 505590 434260
rect 505016 434136 505050 434170
rect 505106 434136 505140 434170
rect 505196 434136 505230 434170
rect 505286 434136 505320 434170
rect 505376 434136 505410 434170
rect 505466 434136 505500 434170
rect 505556 434136 505590 434170
rect 505016 434046 505050 434080
rect 505106 434046 505140 434080
rect 505196 434046 505230 434080
rect 505286 434046 505320 434080
rect 505376 434046 505410 434080
rect 505466 434046 505500 434080
rect 505556 434046 505590 434080
rect 505016 433956 505050 433990
rect 505106 433956 505140 433990
rect 505196 433956 505230 433990
rect 505286 433956 505320 433990
rect 505376 433956 505410 433990
rect 505466 433956 505500 433990
rect 505556 433956 505590 433990
rect 505016 433866 505050 433900
rect 505106 433866 505140 433900
rect 505196 433866 505230 433900
rect 505286 433866 505320 433900
rect 505376 433866 505410 433900
rect 505466 433866 505500 433900
rect 505556 433866 505590 433900
rect 505016 433776 505050 433810
rect 505106 433776 505140 433810
rect 505196 433776 505230 433810
rect 505286 433776 505320 433810
rect 505376 433776 505410 433810
rect 505466 433776 505500 433810
rect 505556 433776 505590 433810
rect 505016 433686 505050 433720
rect 505106 433686 505140 433720
rect 505196 433686 505230 433720
rect 505286 433686 505320 433720
rect 505376 433686 505410 433720
rect 505466 433686 505500 433720
rect 505556 433686 505590 433720
rect 506304 434226 506338 434260
rect 506394 434226 506428 434260
rect 506484 434226 506518 434260
rect 506574 434226 506608 434260
rect 506664 434226 506698 434260
rect 506754 434226 506788 434260
rect 506844 434226 506878 434260
rect 506304 434136 506338 434170
rect 506394 434136 506428 434170
rect 506484 434136 506518 434170
rect 506574 434136 506608 434170
rect 506664 434136 506698 434170
rect 506754 434136 506788 434170
rect 506844 434136 506878 434170
rect 506304 434046 506338 434080
rect 506394 434046 506428 434080
rect 506484 434046 506518 434080
rect 506574 434046 506608 434080
rect 506664 434046 506698 434080
rect 506754 434046 506788 434080
rect 506844 434046 506878 434080
rect 506304 433956 506338 433990
rect 506394 433956 506428 433990
rect 506484 433956 506518 433990
rect 506574 433956 506608 433990
rect 506664 433956 506698 433990
rect 506754 433956 506788 433990
rect 506844 433956 506878 433990
rect 506304 433866 506338 433900
rect 506394 433866 506428 433900
rect 506484 433866 506518 433900
rect 506574 433866 506608 433900
rect 506664 433866 506698 433900
rect 506754 433866 506788 433900
rect 506844 433866 506878 433900
rect 506304 433776 506338 433810
rect 506394 433776 506428 433810
rect 506484 433776 506518 433810
rect 506574 433776 506608 433810
rect 506664 433776 506698 433810
rect 506754 433776 506788 433810
rect 506844 433776 506878 433810
rect 506304 433686 506338 433720
rect 506394 433686 506428 433720
rect 506484 433686 506518 433720
rect 506574 433686 506608 433720
rect 506664 433686 506698 433720
rect 506754 433686 506788 433720
rect 506844 433686 506878 433720
rect 507592 434226 507626 434260
rect 507682 434226 507716 434260
rect 507772 434226 507806 434260
rect 507862 434226 507896 434260
rect 507952 434226 507986 434260
rect 508042 434226 508076 434260
rect 508132 434226 508166 434260
rect 507592 434136 507626 434170
rect 507682 434136 507716 434170
rect 507772 434136 507806 434170
rect 507862 434136 507896 434170
rect 507952 434136 507986 434170
rect 508042 434136 508076 434170
rect 508132 434136 508166 434170
rect 507592 434046 507626 434080
rect 507682 434046 507716 434080
rect 507772 434046 507806 434080
rect 507862 434046 507896 434080
rect 507952 434046 507986 434080
rect 508042 434046 508076 434080
rect 508132 434046 508166 434080
rect 507592 433956 507626 433990
rect 507682 433956 507716 433990
rect 507772 433956 507806 433990
rect 507862 433956 507896 433990
rect 507952 433956 507986 433990
rect 508042 433956 508076 433990
rect 508132 433956 508166 433990
rect 507592 433866 507626 433900
rect 507682 433866 507716 433900
rect 507772 433866 507806 433900
rect 507862 433866 507896 433900
rect 507952 433866 507986 433900
rect 508042 433866 508076 433900
rect 508132 433866 508166 433900
rect 507592 433776 507626 433810
rect 507682 433776 507716 433810
rect 507772 433776 507806 433810
rect 507862 433776 507896 433810
rect 507952 433776 507986 433810
rect 508042 433776 508076 433810
rect 508132 433776 508166 433810
rect 507592 433686 507626 433720
rect 507682 433686 507716 433720
rect 507772 433686 507806 433720
rect 507862 433686 507896 433720
rect 507952 433686 507986 433720
rect 508042 433686 508076 433720
rect 508132 433686 508166 433720
rect 508880 434226 508914 434260
rect 508970 434226 509004 434260
rect 509060 434226 509094 434260
rect 509150 434226 509184 434260
rect 509240 434226 509274 434260
rect 509330 434226 509364 434260
rect 509420 434226 509454 434260
rect 508880 434136 508914 434170
rect 508970 434136 509004 434170
rect 509060 434136 509094 434170
rect 509150 434136 509184 434170
rect 509240 434136 509274 434170
rect 509330 434136 509364 434170
rect 509420 434136 509454 434170
rect 508880 434046 508914 434080
rect 508970 434046 509004 434080
rect 509060 434046 509094 434080
rect 509150 434046 509184 434080
rect 509240 434046 509274 434080
rect 509330 434046 509364 434080
rect 509420 434046 509454 434080
rect 508880 433956 508914 433990
rect 508970 433956 509004 433990
rect 509060 433956 509094 433990
rect 509150 433956 509184 433990
rect 509240 433956 509274 433990
rect 509330 433956 509364 433990
rect 509420 433956 509454 433990
rect 508880 433866 508914 433900
rect 508970 433866 509004 433900
rect 509060 433866 509094 433900
rect 509150 433866 509184 433900
rect 509240 433866 509274 433900
rect 509330 433866 509364 433900
rect 509420 433866 509454 433900
rect 508880 433776 508914 433810
rect 508970 433776 509004 433810
rect 509060 433776 509094 433810
rect 509150 433776 509184 433810
rect 509240 433776 509274 433810
rect 509330 433776 509364 433810
rect 509420 433776 509454 433810
rect 508880 433686 508914 433720
rect 508970 433686 509004 433720
rect 509060 433686 509094 433720
rect 509150 433686 509184 433720
rect 509240 433686 509274 433720
rect 509330 433686 509364 433720
rect 509420 433686 509454 433720
rect 510168 434226 510202 434260
rect 510258 434226 510292 434260
rect 510348 434226 510382 434260
rect 510438 434226 510472 434260
rect 510528 434226 510562 434260
rect 510618 434226 510652 434260
rect 510708 434226 510742 434260
rect 510168 434136 510202 434170
rect 510258 434136 510292 434170
rect 510348 434136 510382 434170
rect 510438 434136 510472 434170
rect 510528 434136 510562 434170
rect 510618 434136 510652 434170
rect 510708 434136 510742 434170
rect 510168 434046 510202 434080
rect 510258 434046 510292 434080
rect 510348 434046 510382 434080
rect 510438 434046 510472 434080
rect 510528 434046 510562 434080
rect 510618 434046 510652 434080
rect 510708 434046 510742 434080
rect 510168 433956 510202 433990
rect 510258 433956 510292 433990
rect 510348 433956 510382 433990
rect 510438 433956 510472 433990
rect 510528 433956 510562 433990
rect 510618 433956 510652 433990
rect 510708 433956 510742 433990
rect 510168 433866 510202 433900
rect 510258 433866 510292 433900
rect 510348 433866 510382 433900
rect 510438 433866 510472 433900
rect 510528 433866 510562 433900
rect 510618 433866 510652 433900
rect 510708 433866 510742 433900
rect 510168 433776 510202 433810
rect 510258 433776 510292 433810
rect 510348 433776 510382 433810
rect 510438 433776 510472 433810
rect 510528 433776 510562 433810
rect 510618 433776 510652 433810
rect 510708 433776 510742 433810
rect 510168 433686 510202 433720
rect 510258 433686 510292 433720
rect 510348 433686 510382 433720
rect 510438 433686 510472 433720
rect 510528 433686 510562 433720
rect 510618 433686 510652 433720
rect 510708 433686 510742 433720
rect 511456 434226 511490 434260
rect 511546 434226 511580 434260
rect 511636 434226 511670 434260
rect 511726 434226 511760 434260
rect 511816 434226 511850 434260
rect 511906 434226 511940 434260
rect 511996 434226 512030 434260
rect 511456 434136 511490 434170
rect 511546 434136 511580 434170
rect 511636 434136 511670 434170
rect 511726 434136 511760 434170
rect 511816 434136 511850 434170
rect 511906 434136 511940 434170
rect 511996 434136 512030 434170
rect 511456 434046 511490 434080
rect 511546 434046 511580 434080
rect 511636 434046 511670 434080
rect 511726 434046 511760 434080
rect 511816 434046 511850 434080
rect 511906 434046 511940 434080
rect 511996 434046 512030 434080
rect 511456 433956 511490 433990
rect 511546 433956 511580 433990
rect 511636 433956 511670 433990
rect 511726 433956 511760 433990
rect 511816 433956 511850 433990
rect 511906 433956 511940 433990
rect 511996 433956 512030 433990
rect 511456 433866 511490 433900
rect 511546 433866 511580 433900
rect 511636 433866 511670 433900
rect 511726 433866 511760 433900
rect 511816 433866 511850 433900
rect 511906 433866 511940 433900
rect 511996 433866 512030 433900
rect 511456 433776 511490 433810
rect 511546 433776 511580 433810
rect 511636 433776 511670 433810
rect 511726 433776 511760 433810
rect 511816 433776 511850 433810
rect 511906 433776 511940 433810
rect 511996 433776 512030 433810
rect 511456 433686 511490 433720
rect 511546 433686 511580 433720
rect 511636 433686 511670 433720
rect 511726 433686 511760 433720
rect 511816 433686 511850 433720
rect 511906 433686 511940 433720
rect 511996 433686 512030 433720
rect 512744 434226 512778 434260
rect 512834 434226 512868 434260
rect 512924 434226 512958 434260
rect 513014 434226 513048 434260
rect 513104 434226 513138 434260
rect 513194 434226 513228 434260
rect 513284 434226 513318 434260
rect 512744 434136 512778 434170
rect 512834 434136 512868 434170
rect 512924 434136 512958 434170
rect 513014 434136 513048 434170
rect 513104 434136 513138 434170
rect 513194 434136 513228 434170
rect 513284 434136 513318 434170
rect 512744 434046 512778 434080
rect 512834 434046 512868 434080
rect 512924 434046 512958 434080
rect 513014 434046 513048 434080
rect 513104 434046 513138 434080
rect 513194 434046 513228 434080
rect 513284 434046 513318 434080
rect 512744 433956 512778 433990
rect 512834 433956 512868 433990
rect 512924 433956 512958 433990
rect 513014 433956 513048 433990
rect 513104 433956 513138 433990
rect 513194 433956 513228 433990
rect 513284 433956 513318 433990
rect 512744 433866 512778 433900
rect 512834 433866 512868 433900
rect 512924 433866 512958 433900
rect 513014 433866 513048 433900
rect 513104 433866 513138 433900
rect 513194 433866 513228 433900
rect 513284 433866 513318 433900
rect 512744 433776 512778 433810
rect 512834 433776 512868 433810
rect 512924 433776 512958 433810
rect 513014 433776 513048 433810
rect 513104 433776 513138 433810
rect 513194 433776 513228 433810
rect 513284 433776 513318 433810
rect 512744 433686 512778 433720
rect 512834 433686 512868 433720
rect 512924 433686 512958 433720
rect 513014 433686 513048 433720
rect 513104 433686 513138 433720
rect 513194 433686 513228 433720
rect 513284 433686 513318 433720
rect 503728 432938 503762 432972
rect 503818 432938 503852 432972
rect 503908 432938 503942 432972
rect 503998 432938 504032 432972
rect 504088 432938 504122 432972
rect 504178 432938 504212 432972
rect 504268 432938 504302 432972
rect 503728 432848 503762 432882
rect 503818 432848 503852 432882
rect 503908 432848 503942 432882
rect 503998 432848 504032 432882
rect 504088 432848 504122 432882
rect 504178 432848 504212 432882
rect 504268 432848 504302 432882
rect 503728 432758 503762 432792
rect 503818 432758 503852 432792
rect 503908 432758 503942 432792
rect 503998 432758 504032 432792
rect 504088 432758 504122 432792
rect 504178 432758 504212 432792
rect 504268 432758 504302 432792
rect 503728 432668 503762 432702
rect 503818 432668 503852 432702
rect 503908 432668 503942 432702
rect 503998 432668 504032 432702
rect 504088 432668 504122 432702
rect 504178 432668 504212 432702
rect 504268 432668 504302 432702
rect 503728 432578 503762 432612
rect 503818 432578 503852 432612
rect 503908 432578 503942 432612
rect 503998 432578 504032 432612
rect 504088 432578 504122 432612
rect 504178 432578 504212 432612
rect 504268 432578 504302 432612
rect 503728 432488 503762 432522
rect 503818 432488 503852 432522
rect 503908 432488 503942 432522
rect 503998 432488 504032 432522
rect 504088 432488 504122 432522
rect 504178 432488 504212 432522
rect 504268 432488 504302 432522
rect 503728 432398 503762 432432
rect 503818 432398 503852 432432
rect 503908 432398 503942 432432
rect 503998 432398 504032 432432
rect 504088 432398 504122 432432
rect 504178 432398 504212 432432
rect 504268 432398 504302 432432
rect 505016 432938 505050 432972
rect 505106 432938 505140 432972
rect 505196 432938 505230 432972
rect 505286 432938 505320 432972
rect 505376 432938 505410 432972
rect 505466 432938 505500 432972
rect 505556 432938 505590 432972
rect 505016 432848 505050 432882
rect 505106 432848 505140 432882
rect 505196 432848 505230 432882
rect 505286 432848 505320 432882
rect 505376 432848 505410 432882
rect 505466 432848 505500 432882
rect 505556 432848 505590 432882
rect 505016 432758 505050 432792
rect 505106 432758 505140 432792
rect 505196 432758 505230 432792
rect 505286 432758 505320 432792
rect 505376 432758 505410 432792
rect 505466 432758 505500 432792
rect 505556 432758 505590 432792
rect 505016 432668 505050 432702
rect 505106 432668 505140 432702
rect 505196 432668 505230 432702
rect 505286 432668 505320 432702
rect 505376 432668 505410 432702
rect 505466 432668 505500 432702
rect 505556 432668 505590 432702
rect 505016 432578 505050 432612
rect 505106 432578 505140 432612
rect 505196 432578 505230 432612
rect 505286 432578 505320 432612
rect 505376 432578 505410 432612
rect 505466 432578 505500 432612
rect 505556 432578 505590 432612
rect 505016 432488 505050 432522
rect 505106 432488 505140 432522
rect 505196 432488 505230 432522
rect 505286 432488 505320 432522
rect 505376 432488 505410 432522
rect 505466 432488 505500 432522
rect 505556 432488 505590 432522
rect 505016 432398 505050 432432
rect 505106 432398 505140 432432
rect 505196 432398 505230 432432
rect 505286 432398 505320 432432
rect 505376 432398 505410 432432
rect 505466 432398 505500 432432
rect 505556 432398 505590 432432
rect 506304 432938 506338 432972
rect 506394 432938 506428 432972
rect 506484 432938 506518 432972
rect 506574 432938 506608 432972
rect 506664 432938 506698 432972
rect 506754 432938 506788 432972
rect 506844 432938 506878 432972
rect 506304 432848 506338 432882
rect 506394 432848 506428 432882
rect 506484 432848 506518 432882
rect 506574 432848 506608 432882
rect 506664 432848 506698 432882
rect 506754 432848 506788 432882
rect 506844 432848 506878 432882
rect 506304 432758 506338 432792
rect 506394 432758 506428 432792
rect 506484 432758 506518 432792
rect 506574 432758 506608 432792
rect 506664 432758 506698 432792
rect 506754 432758 506788 432792
rect 506844 432758 506878 432792
rect 506304 432668 506338 432702
rect 506394 432668 506428 432702
rect 506484 432668 506518 432702
rect 506574 432668 506608 432702
rect 506664 432668 506698 432702
rect 506754 432668 506788 432702
rect 506844 432668 506878 432702
rect 506304 432578 506338 432612
rect 506394 432578 506428 432612
rect 506484 432578 506518 432612
rect 506574 432578 506608 432612
rect 506664 432578 506698 432612
rect 506754 432578 506788 432612
rect 506844 432578 506878 432612
rect 506304 432488 506338 432522
rect 506394 432488 506428 432522
rect 506484 432488 506518 432522
rect 506574 432488 506608 432522
rect 506664 432488 506698 432522
rect 506754 432488 506788 432522
rect 506844 432488 506878 432522
rect 506304 432398 506338 432432
rect 506394 432398 506428 432432
rect 506484 432398 506518 432432
rect 506574 432398 506608 432432
rect 506664 432398 506698 432432
rect 506754 432398 506788 432432
rect 506844 432398 506878 432432
rect 507592 432938 507626 432972
rect 507682 432938 507716 432972
rect 507772 432938 507806 432972
rect 507862 432938 507896 432972
rect 507952 432938 507986 432972
rect 508042 432938 508076 432972
rect 508132 432938 508166 432972
rect 507592 432848 507626 432882
rect 507682 432848 507716 432882
rect 507772 432848 507806 432882
rect 507862 432848 507896 432882
rect 507952 432848 507986 432882
rect 508042 432848 508076 432882
rect 508132 432848 508166 432882
rect 507592 432758 507626 432792
rect 507682 432758 507716 432792
rect 507772 432758 507806 432792
rect 507862 432758 507896 432792
rect 507952 432758 507986 432792
rect 508042 432758 508076 432792
rect 508132 432758 508166 432792
rect 507592 432668 507626 432702
rect 507682 432668 507716 432702
rect 507772 432668 507806 432702
rect 507862 432668 507896 432702
rect 507952 432668 507986 432702
rect 508042 432668 508076 432702
rect 508132 432668 508166 432702
rect 507592 432578 507626 432612
rect 507682 432578 507716 432612
rect 507772 432578 507806 432612
rect 507862 432578 507896 432612
rect 507952 432578 507986 432612
rect 508042 432578 508076 432612
rect 508132 432578 508166 432612
rect 507592 432488 507626 432522
rect 507682 432488 507716 432522
rect 507772 432488 507806 432522
rect 507862 432488 507896 432522
rect 507952 432488 507986 432522
rect 508042 432488 508076 432522
rect 508132 432488 508166 432522
rect 507592 432398 507626 432432
rect 507682 432398 507716 432432
rect 507772 432398 507806 432432
rect 507862 432398 507896 432432
rect 507952 432398 507986 432432
rect 508042 432398 508076 432432
rect 508132 432398 508166 432432
rect 508880 432938 508914 432972
rect 508970 432938 509004 432972
rect 509060 432938 509094 432972
rect 509150 432938 509184 432972
rect 509240 432938 509274 432972
rect 509330 432938 509364 432972
rect 509420 432938 509454 432972
rect 508880 432848 508914 432882
rect 508970 432848 509004 432882
rect 509060 432848 509094 432882
rect 509150 432848 509184 432882
rect 509240 432848 509274 432882
rect 509330 432848 509364 432882
rect 509420 432848 509454 432882
rect 508880 432758 508914 432792
rect 508970 432758 509004 432792
rect 509060 432758 509094 432792
rect 509150 432758 509184 432792
rect 509240 432758 509274 432792
rect 509330 432758 509364 432792
rect 509420 432758 509454 432792
rect 508880 432668 508914 432702
rect 508970 432668 509004 432702
rect 509060 432668 509094 432702
rect 509150 432668 509184 432702
rect 509240 432668 509274 432702
rect 509330 432668 509364 432702
rect 509420 432668 509454 432702
rect 508880 432578 508914 432612
rect 508970 432578 509004 432612
rect 509060 432578 509094 432612
rect 509150 432578 509184 432612
rect 509240 432578 509274 432612
rect 509330 432578 509364 432612
rect 509420 432578 509454 432612
rect 508880 432488 508914 432522
rect 508970 432488 509004 432522
rect 509060 432488 509094 432522
rect 509150 432488 509184 432522
rect 509240 432488 509274 432522
rect 509330 432488 509364 432522
rect 509420 432488 509454 432522
rect 508880 432398 508914 432432
rect 508970 432398 509004 432432
rect 509060 432398 509094 432432
rect 509150 432398 509184 432432
rect 509240 432398 509274 432432
rect 509330 432398 509364 432432
rect 509420 432398 509454 432432
rect 510168 432938 510202 432972
rect 510258 432938 510292 432972
rect 510348 432938 510382 432972
rect 510438 432938 510472 432972
rect 510528 432938 510562 432972
rect 510618 432938 510652 432972
rect 510708 432938 510742 432972
rect 510168 432848 510202 432882
rect 510258 432848 510292 432882
rect 510348 432848 510382 432882
rect 510438 432848 510472 432882
rect 510528 432848 510562 432882
rect 510618 432848 510652 432882
rect 510708 432848 510742 432882
rect 510168 432758 510202 432792
rect 510258 432758 510292 432792
rect 510348 432758 510382 432792
rect 510438 432758 510472 432792
rect 510528 432758 510562 432792
rect 510618 432758 510652 432792
rect 510708 432758 510742 432792
rect 510168 432668 510202 432702
rect 510258 432668 510292 432702
rect 510348 432668 510382 432702
rect 510438 432668 510472 432702
rect 510528 432668 510562 432702
rect 510618 432668 510652 432702
rect 510708 432668 510742 432702
rect 510168 432578 510202 432612
rect 510258 432578 510292 432612
rect 510348 432578 510382 432612
rect 510438 432578 510472 432612
rect 510528 432578 510562 432612
rect 510618 432578 510652 432612
rect 510708 432578 510742 432612
rect 510168 432488 510202 432522
rect 510258 432488 510292 432522
rect 510348 432488 510382 432522
rect 510438 432488 510472 432522
rect 510528 432488 510562 432522
rect 510618 432488 510652 432522
rect 510708 432488 510742 432522
rect 510168 432398 510202 432432
rect 510258 432398 510292 432432
rect 510348 432398 510382 432432
rect 510438 432398 510472 432432
rect 510528 432398 510562 432432
rect 510618 432398 510652 432432
rect 510708 432398 510742 432432
rect 511456 432938 511490 432972
rect 511546 432938 511580 432972
rect 511636 432938 511670 432972
rect 511726 432938 511760 432972
rect 511816 432938 511850 432972
rect 511906 432938 511940 432972
rect 511996 432938 512030 432972
rect 511456 432848 511490 432882
rect 511546 432848 511580 432882
rect 511636 432848 511670 432882
rect 511726 432848 511760 432882
rect 511816 432848 511850 432882
rect 511906 432848 511940 432882
rect 511996 432848 512030 432882
rect 511456 432758 511490 432792
rect 511546 432758 511580 432792
rect 511636 432758 511670 432792
rect 511726 432758 511760 432792
rect 511816 432758 511850 432792
rect 511906 432758 511940 432792
rect 511996 432758 512030 432792
rect 511456 432668 511490 432702
rect 511546 432668 511580 432702
rect 511636 432668 511670 432702
rect 511726 432668 511760 432702
rect 511816 432668 511850 432702
rect 511906 432668 511940 432702
rect 511996 432668 512030 432702
rect 511456 432578 511490 432612
rect 511546 432578 511580 432612
rect 511636 432578 511670 432612
rect 511726 432578 511760 432612
rect 511816 432578 511850 432612
rect 511906 432578 511940 432612
rect 511996 432578 512030 432612
rect 511456 432488 511490 432522
rect 511546 432488 511580 432522
rect 511636 432488 511670 432522
rect 511726 432488 511760 432522
rect 511816 432488 511850 432522
rect 511906 432488 511940 432522
rect 511996 432488 512030 432522
rect 511456 432398 511490 432432
rect 511546 432398 511580 432432
rect 511636 432398 511670 432432
rect 511726 432398 511760 432432
rect 511816 432398 511850 432432
rect 511906 432398 511940 432432
rect 511996 432398 512030 432432
rect 512744 432938 512778 432972
rect 512834 432938 512868 432972
rect 512924 432938 512958 432972
rect 513014 432938 513048 432972
rect 513104 432938 513138 432972
rect 513194 432938 513228 432972
rect 513284 432938 513318 432972
rect 512744 432848 512778 432882
rect 512834 432848 512868 432882
rect 512924 432848 512958 432882
rect 513014 432848 513048 432882
rect 513104 432848 513138 432882
rect 513194 432848 513228 432882
rect 513284 432848 513318 432882
rect 512744 432758 512778 432792
rect 512834 432758 512868 432792
rect 512924 432758 512958 432792
rect 513014 432758 513048 432792
rect 513104 432758 513138 432792
rect 513194 432758 513228 432792
rect 513284 432758 513318 432792
rect 512744 432668 512778 432702
rect 512834 432668 512868 432702
rect 512924 432668 512958 432702
rect 513014 432668 513048 432702
rect 513104 432668 513138 432702
rect 513194 432668 513228 432702
rect 513284 432668 513318 432702
rect 512744 432578 512778 432612
rect 512834 432578 512868 432612
rect 512924 432578 512958 432612
rect 513014 432578 513048 432612
rect 513104 432578 513138 432612
rect 513194 432578 513228 432612
rect 513284 432578 513318 432612
rect 512744 432488 512778 432522
rect 512834 432488 512868 432522
rect 512924 432488 512958 432522
rect 513014 432488 513048 432522
rect 513104 432488 513138 432522
rect 513194 432488 513228 432522
rect 513284 432488 513318 432522
rect 512744 432398 512778 432432
rect 512834 432398 512868 432432
rect 512924 432398 512958 432432
rect 513014 432398 513048 432432
rect 513104 432398 513138 432432
rect 513194 432398 513228 432432
rect 513284 432398 513318 432432
rect 562270 454112 562304 455088
rect 562528 454112 562562 455088
rect 562786 454112 562820 455088
rect 563044 454112 563078 455088
rect 563302 454112 563336 455088
rect 563560 454112 563594 455088
rect 563818 454112 563852 455088
rect 564076 454112 564110 455088
rect 564334 454112 564368 455088
rect 564592 454112 564626 455088
rect 564850 454112 564884 455088
rect 565108 454112 565142 455088
rect 565366 454112 565400 455088
rect 565624 454112 565658 455088
rect 565882 454112 565916 455088
rect 566140 454112 566174 455088
rect 566398 454112 566432 455088
rect 566656 454112 566690 455088
rect 566914 454112 566948 455088
rect 567172 454112 567206 455088
rect 567430 454112 567464 455088
<< psubdiff >>
rect 572316 495514 572412 495548
rect 577642 495514 577738 495548
rect 572316 495452 572350 495514
rect 577704 495452 577738 495514
rect 572316 494296 572350 494358
rect 577704 494296 577738 494358
rect 572316 494262 572412 494296
rect 577642 494262 577738 494296
rect 527568 475332 528616 475356
rect 500344 475308 501392 475332
rect 500344 432068 500368 475308
rect 501368 432068 501392 475308
rect 502368 475284 526568 475308
rect 502368 474284 502392 475284
rect 526544 474284 526568 475284
rect 502368 474260 526568 474284
rect 507162 473280 507286 473284
rect 506508 473256 507286 473280
rect 506508 472856 506532 473256
rect 507108 472856 507286 473256
rect 506508 472832 507286 472856
rect 507162 471870 507286 472832
rect 507162 470878 507186 471870
rect 507262 470878 507286 471870
rect 507162 469914 507286 470878
rect 506508 469890 507286 469914
rect 506508 469490 506532 469890
rect 507108 469490 507286 469890
rect 506508 469466 507286 469490
rect 507162 469464 507286 469466
rect 525672 472468 526486 472492
rect 510452 468834 510832 468858
rect 506368 468386 508168 468436
rect 506368 468286 506468 468386
rect 508068 468286 508168 468386
rect 506368 468236 508168 468286
rect 506368 462886 508168 462936
rect 506368 462786 506468 462886
rect 508068 462786 508168 462886
rect 506368 462736 508168 462786
rect 510452 462382 510476 468834
rect 510808 462382 510832 468834
rect 510452 462358 510832 462382
rect 525672 461284 525696 472468
rect 526462 461284 526486 472468
rect 525672 461260 526486 461284
rect 516598 460708 522950 460732
rect 516598 460138 516622 460708
rect 522926 460138 522950 460708
rect 516598 460114 522950 460138
rect 516598 457464 522950 457488
rect 516598 456894 516622 457464
rect 522926 456894 522950 457464
rect 516598 456870 522950 456894
rect 516598 452504 522950 452528
rect 516598 451934 516622 452504
rect 522926 451934 522950 452504
rect 516598 451910 522950 451934
rect 500344 432044 501392 432068
rect 503370 438448 513674 438482
rect 503370 438414 503486 438448
rect 503520 438414 503576 438448
rect 503610 438414 503666 438448
rect 503700 438414 503756 438448
rect 503790 438414 503846 438448
rect 503880 438414 503936 438448
rect 503970 438414 504026 438448
rect 504060 438414 504116 438448
rect 504150 438414 504206 438448
rect 504240 438414 504296 438448
rect 504330 438414 504386 438448
rect 504420 438414 504476 438448
rect 504510 438414 504566 438448
rect 504600 438414 504774 438448
rect 504808 438414 504864 438448
rect 504898 438414 504954 438448
rect 504988 438414 505044 438448
rect 505078 438414 505134 438448
rect 505168 438414 505224 438448
rect 505258 438414 505314 438448
rect 505348 438414 505404 438448
rect 505438 438414 505494 438448
rect 505528 438414 505584 438448
rect 505618 438414 505674 438448
rect 505708 438414 505764 438448
rect 505798 438414 505854 438448
rect 505888 438414 506062 438448
rect 506096 438414 506152 438448
rect 506186 438414 506242 438448
rect 506276 438414 506332 438448
rect 506366 438414 506422 438448
rect 506456 438414 506512 438448
rect 506546 438414 506602 438448
rect 506636 438414 506692 438448
rect 506726 438414 506782 438448
rect 506816 438414 506872 438448
rect 506906 438414 506962 438448
rect 506996 438414 507052 438448
rect 507086 438414 507142 438448
rect 507176 438414 507350 438448
rect 507384 438414 507440 438448
rect 507474 438414 507530 438448
rect 507564 438414 507620 438448
rect 507654 438414 507710 438448
rect 507744 438414 507800 438448
rect 507834 438414 507890 438448
rect 507924 438414 507980 438448
rect 508014 438414 508070 438448
rect 508104 438414 508160 438448
rect 508194 438414 508250 438448
rect 508284 438414 508340 438448
rect 508374 438414 508430 438448
rect 508464 438414 508638 438448
rect 508672 438414 508728 438448
rect 508762 438414 508818 438448
rect 508852 438414 508908 438448
rect 508942 438414 508998 438448
rect 509032 438414 509088 438448
rect 509122 438414 509178 438448
rect 509212 438414 509268 438448
rect 509302 438414 509358 438448
rect 509392 438414 509448 438448
rect 509482 438414 509538 438448
rect 509572 438414 509628 438448
rect 509662 438414 509718 438448
rect 509752 438414 509926 438448
rect 509960 438414 510016 438448
rect 510050 438414 510106 438448
rect 510140 438414 510196 438448
rect 510230 438414 510286 438448
rect 510320 438414 510376 438448
rect 510410 438414 510466 438448
rect 510500 438414 510556 438448
rect 510590 438414 510646 438448
rect 510680 438414 510736 438448
rect 510770 438414 510826 438448
rect 510860 438414 510916 438448
rect 510950 438414 511006 438448
rect 511040 438414 511214 438448
rect 511248 438414 511304 438448
rect 511338 438414 511394 438448
rect 511428 438414 511484 438448
rect 511518 438414 511574 438448
rect 511608 438414 511664 438448
rect 511698 438414 511754 438448
rect 511788 438414 511844 438448
rect 511878 438414 511934 438448
rect 511968 438414 512024 438448
rect 512058 438414 512114 438448
rect 512148 438414 512204 438448
rect 512238 438414 512294 438448
rect 512328 438414 512502 438448
rect 512536 438414 512592 438448
rect 512626 438414 512682 438448
rect 512716 438414 512772 438448
rect 512806 438414 512862 438448
rect 512896 438414 512952 438448
rect 512986 438414 513042 438448
rect 513076 438414 513132 438448
rect 513166 438414 513222 438448
rect 513256 438414 513312 438448
rect 513346 438414 513402 438448
rect 513436 438414 513492 438448
rect 513526 438414 513582 438448
rect 513616 438414 513674 438448
rect 503370 438381 513674 438414
rect 503370 438352 503471 438381
rect 503370 438318 503402 438352
rect 503436 438318 503471 438352
rect 504557 438352 504759 438381
rect 503370 438262 503471 438318
rect 503370 438228 503402 438262
rect 503436 438228 503471 438262
rect 503370 438172 503471 438228
rect 503370 438138 503402 438172
rect 503436 438138 503471 438172
rect 503370 438082 503471 438138
rect 503370 438048 503402 438082
rect 503436 438048 503471 438082
rect 503370 437992 503471 438048
rect 503370 437958 503402 437992
rect 503436 437958 503471 437992
rect 503370 437902 503471 437958
rect 503370 437868 503402 437902
rect 503436 437868 503471 437902
rect 503370 437812 503471 437868
rect 503370 437778 503402 437812
rect 503436 437778 503471 437812
rect 503370 437722 503471 437778
rect 503370 437688 503402 437722
rect 503436 437688 503471 437722
rect 503370 437632 503471 437688
rect 503370 437598 503402 437632
rect 503436 437598 503471 437632
rect 503370 437542 503471 437598
rect 503370 437508 503402 437542
rect 503436 437508 503471 437542
rect 503370 437452 503471 437508
rect 503370 437418 503402 437452
rect 503436 437418 503471 437452
rect 503370 437362 503471 437418
rect 503370 437328 503402 437362
rect 503436 437328 503471 437362
rect 504557 438318 504589 438352
rect 504623 438318 504690 438352
rect 504724 438318 504759 438352
rect 505845 438352 506047 438381
rect 504557 438262 504759 438318
rect 504557 438228 504589 438262
rect 504623 438228 504690 438262
rect 504724 438228 504759 438262
rect 504557 438172 504759 438228
rect 504557 438138 504589 438172
rect 504623 438138 504690 438172
rect 504724 438138 504759 438172
rect 504557 438082 504759 438138
rect 504557 438048 504589 438082
rect 504623 438048 504690 438082
rect 504724 438048 504759 438082
rect 504557 437992 504759 438048
rect 504557 437958 504589 437992
rect 504623 437958 504690 437992
rect 504724 437958 504759 437992
rect 504557 437902 504759 437958
rect 504557 437868 504589 437902
rect 504623 437868 504690 437902
rect 504724 437868 504759 437902
rect 504557 437812 504759 437868
rect 504557 437778 504589 437812
rect 504623 437778 504690 437812
rect 504724 437778 504759 437812
rect 504557 437722 504759 437778
rect 504557 437688 504589 437722
rect 504623 437688 504690 437722
rect 504724 437688 504759 437722
rect 504557 437632 504759 437688
rect 504557 437598 504589 437632
rect 504623 437598 504690 437632
rect 504724 437598 504759 437632
rect 504557 437542 504759 437598
rect 504557 437508 504589 437542
rect 504623 437508 504690 437542
rect 504724 437508 504759 437542
rect 504557 437452 504759 437508
rect 504557 437418 504589 437452
rect 504623 437418 504690 437452
rect 504724 437418 504759 437452
rect 504557 437362 504759 437418
rect 503370 437295 503471 437328
rect 504557 437328 504589 437362
rect 504623 437328 504690 437362
rect 504724 437328 504759 437362
rect 505845 438318 505877 438352
rect 505911 438318 505978 438352
rect 506012 438318 506047 438352
rect 507133 438352 507335 438381
rect 505845 438262 506047 438318
rect 505845 438228 505877 438262
rect 505911 438228 505978 438262
rect 506012 438228 506047 438262
rect 505845 438172 506047 438228
rect 505845 438138 505877 438172
rect 505911 438138 505978 438172
rect 506012 438138 506047 438172
rect 505845 438082 506047 438138
rect 505845 438048 505877 438082
rect 505911 438048 505978 438082
rect 506012 438048 506047 438082
rect 505845 437992 506047 438048
rect 505845 437958 505877 437992
rect 505911 437958 505978 437992
rect 506012 437958 506047 437992
rect 505845 437902 506047 437958
rect 505845 437868 505877 437902
rect 505911 437868 505978 437902
rect 506012 437868 506047 437902
rect 505845 437812 506047 437868
rect 505845 437778 505877 437812
rect 505911 437778 505978 437812
rect 506012 437778 506047 437812
rect 505845 437722 506047 437778
rect 505845 437688 505877 437722
rect 505911 437688 505978 437722
rect 506012 437688 506047 437722
rect 505845 437632 506047 437688
rect 505845 437598 505877 437632
rect 505911 437598 505978 437632
rect 506012 437598 506047 437632
rect 505845 437542 506047 437598
rect 505845 437508 505877 437542
rect 505911 437508 505978 437542
rect 506012 437508 506047 437542
rect 505845 437452 506047 437508
rect 505845 437418 505877 437452
rect 505911 437418 505978 437452
rect 506012 437418 506047 437452
rect 505845 437362 506047 437418
rect 504557 437295 504759 437328
rect 505845 437328 505877 437362
rect 505911 437328 505978 437362
rect 506012 437328 506047 437362
rect 507133 438318 507165 438352
rect 507199 438318 507266 438352
rect 507300 438318 507335 438352
rect 508421 438352 508623 438381
rect 507133 438262 507335 438318
rect 507133 438228 507165 438262
rect 507199 438228 507266 438262
rect 507300 438228 507335 438262
rect 507133 438172 507335 438228
rect 507133 438138 507165 438172
rect 507199 438138 507266 438172
rect 507300 438138 507335 438172
rect 507133 438082 507335 438138
rect 507133 438048 507165 438082
rect 507199 438048 507266 438082
rect 507300 438048 507335 438082
rect 507133 437992 507335 438048
rect 507133 437958 507165 437992
rect 507199 437958 507266 437992
rect 507300 437958 507335 437992
rect 507133 437902 507335 437958
rect 507133 437868 507165 437902
rect 507199 437868 507266 437902
rect 507300 437868 507335 437902
rect 507133 437812 507335 437868
rect 507133 437778 507165 437812
rect 507199 437778 507266 437812
rect 507300 437778 507335 437812
rect 507133 437722 507335 437778
rect 507133 437688 507165 437722
rect 507199 437688 507266 437722
rect 507300 437688 507335 437722
rect 507133 437632 507335 437688
rect 507133 437598 507165 437632
rect 507199 437598 507266 437632
rect 507300 437598 507335 437632
rect 507133 437542 507335 437598
rect 507133 437508 507165 437542
rect 507199 437508 507266 437542
rect 507300 437508 507335 437542
rect 507133 437452 507335 437508
rect 507133 437418 507165 437452
rect 507199 437418 507266 437452
rect 507300 437418 507335 437452
rect 507133 437362 507335 437418
rect 505845 437295 506047 437328
rect 507133 437328 507165 437362
rect 507199 437328 507266 437362
rect 507300 437328 507335 437362
rect 508421 438318 508453 438352
rect 508487 438318 508554 438352
rect 508588 438318 508623 438352
rect 509709 438352 509911 438381
rect 508421 438262 508623 438318
rect 508421 438228 508453 438262
rect 508487 438228 508554 438262
rect 508588 438228 508623 438262
rect 508421 438172 508623 438228
rect 508421 438138 508453 438172
rect 508487 438138 508554 438172
rect 508588 438138 508623 438172
rect 508421 438082 508623 438138
rect 508421 438048 508453 438082
rect 508487 438048 508554 438082
rect 508588 438048 508623 438082
rect 508421 437992 508623 438048
rect 508421 437958 508453 437992
rect 508487 437958 508554 437992
rect 508588 437958 508623 437992
rect 508421 437902 508623 437958
rect 508421 437868 508453 437902
rect 508487 437868 508554 437902
rect 508588 437868 508623 437902
rect 508421 437812 508623 437868
rect 508421 437778 508453 437812
rect 508487 437778 508554 437812
rect 508588 437778 508623 437812
rect 508421 437722 508623 437778
rect 508421 437688 508453 437722
rect 508487 437688 508554 437722
rect 508588 437688 508623 437722
rect 508421 437632 508623 437688
rect 508421 437598 508453 437632
rect 508487 437598 508554 437632
rect 508588 437598 508623 437632
rect 508421 437542 508623 437598
rect 508421 437508 508453 437542
rect 508487 437508 508554 437542
rect 508588 437508 508623 437542
rect 508421 437452 508623 437508
rect 508421 437418 508453 437452
rect 508487 437418 508554 437452
rect 508588 437418 508623 437452
rect 508421 437362 508623 437418
rect 507133 437295 507335 437328
rect 508421 437328 508453 437362
rect 508487 437328 508554 437362
rect 508588 437328 508623 437362
rect 509709 438318 509741 438352
rect 509775 438318 509842 438352
rect 509876 438318 509911 438352
rect 510997 438352 511199 438381
rect 509709 438262 509911 438318
rect 509709 438228 509741 438262
rect 509775 438228 509842 438262
rect 509876 438228 509911 438262
rect 509709 438172 509911 438228
rect 509709 438138 509741 438172
rect 509775 438138 509842 438172
rect 509876 438138 509911 438172
rect 509709 438082 509911 438138
rect 509709 438048 509741 438082
rect 509775 438048 509842 438082
rect 509876 438048 509911 438082
rect 509709 437992 509911 438048
rect 509709 437958 509741 437992
rect 509775 437958 509842 437992
rect 509876 437958 509911 437992
rect 509709 437902 509911 437958
rect 509709 437868 509741 437902
rect 509775 437868 509842 437902
rect 509876 437868 509911 437902
rect 509709 437812 509911 437868
rect 509709 437778 509741 437812
rect 509775 437778 509842 437812
rect 509876 437778 509911 437812
rect 509709 437722 509911 437778
rect 509709 437688 509741 437722
rect 509775 437688 509842 437722
rect 509876 437688 509911 437722
rect 509709 437632 509911 437688
rect 509709 437598 509741 437632
rect 509775 437598 509842 437632
rect 509876 437598 509911 437632
rect 509709 437542 509911 437598
rect 509709 437508 509741 437542
rect 509775 437508 509842 437542
rect 509876 437508 509911 437542
rect 509709 437452 509911 437508
rect 509709 437418 509741 437452
rect 509775 437418 509842 437452
rect 509876 437418 509911 437452
rect 509709 437362 509911 437418
rect 508421 437295 508623 437328
rect 509709 437328 509741 437362
rect 509775 437328 509842 437362
rect 509876 437328 509911 437362
rect 510997 438318 511029 438352
rect 511063 438318 511130 438352
rect 511164 438318 511199 438352
rect 512285 438352 512487 438381
rect 510997 438262 511199 438318
rect 510997 438228 511029 438262
rect 511063 438228 511130 438262
rect 511164 438228 511199 438262
rect 510997 438172 511199 438228
rect 510997 438138 511029 438172
rect 511063 438138 511130 438172
rect 511164 438138 511199 438172
rect 510997 438082 511199 438138
rect 510997 438048 511029 438082
rect 511063 438048 511130 438082
rect 511164 438048 511199 438082
rect 510997 437992 511199 438048
rect 510997 437958 511029 437992
rect 511063 437958 511130 437992
rect 511164 437958 511199 437992
rect 510997 437902 511199 437958
rect 510997 437868 511029 437902
rect 511063 437868 511130 437902
rect 511164 437868 511199 437902
rect 510997 437812 511199 437868
rect 510997 437778 511029 437812
rect 511063 437778 511130 437812
rect 511164 437778 511199 437812
rect 510997 437722 511199 437778
rect 510997 437688 511029 437722
rect 511063 437688 511130 437722
rect 511164 437688 511199 437722
rect 510997 437632 511199 437688
rect 510997 437598 511029 437632
rect 511063 437598 511130 437632
rect 511164 437598 511199 437632
rect 510997 437542 511199 437598
rect 510997 437508 511029 437542
rect 511063 437508 511130 437542
rect 511164 437508 511199 437542
rect 510997 437452 511199 437508
rect 510997 437418 511029 437452
rect 511063 437418 511130 437452
rect 511164 437418 511199 437452
rect 510997 437362 511199 437418
rect 509709 437295 509911 437328
rect 510997 437328 511029 437362
rect 511063 437328 511130 437362
rect 511164 437328 511199 437362
rect 512285 438318 512317 438352
rect 512351 438318 512418 438352
rect 512452 438318 512487 438352
rect 513573 438352 513674 438381
rect 512285 438262 512487 438318
rect 512285 438228 512317 438262
rect 512351 438228 512418 438262
rect 512452 438228 512487 438262
rect 512285 438172 512487 438228
rect 512285 438138 512317 438172
rect 512351 438138 512418 438172
rect 512452 438138 512487 438172
rect 512285 438082 512487 438138
rect 512285 438048 512317 438082
rect 512351 438048 512418 438082
rect 512452 438048 512487 438082
rect 512285 437992 512487 438048
rect 512285 437958 512317 437992
rect 512351 437958 512418 437992
rect 512452 437958 512487 437992
rect 512285 437902 512487 437958
rect 512285 437868 512317 437902
rect 512351 437868 512418 437902
rect 512452 437868 512487 437902
rect 512285 437812 512487 437868
rect 512285 437778 512317 437812
rect 512351 437778 512418 437812
rect 512452 437778 512487 437812
rect 512285 437722 512487 437778
rect 512285 437688 512317 437722
rect 512351 437688 512418 437722
rect 512452 437688 512487 437722
rect 512285 437632 512487 437688
rect 512285 437598 512317 437632
rect 512351 437598 512418 437632
rect 512452 437598 512487 437632
rect 512285 437542 512487 437598
rect 512285 437508 512317 437542
rect 512351 437508 512418 437542
rect 512452 437508 512487 437542
rect 512285 437452 512487 437508
rect 512285 437418 512317 437452
rect 512351 437418 512418 437452
rect 512452 437418 512487 437452
rect 512285 437362 512487 437418
rect 510997 437295 511199 437328
rect 512285 437328 512317 437362
rect 512351 437328 512418 437362
rect 512452 437328 512487 437362
rect 513573 438318 513605 438352
rect 513639 438318 513674 438352
rect 513573 438262 513674 438318
rect 513573 438228 513605 438262
rect 513639 438228 513674 438262
rect 513573 438172 513674 438228
rect 513573 438138 513605 438172
rect 513639 438138 513674 438172
rect 513573 438082 513674 438138
rect 513573 438048 513605 438082
rect 513639 438048 513674 438082
rect 513573 437992 513674 438048
rect 513573 437958 513605 437992
rect 513639 437958 513674 437992
rect 513573 437902 513674 437958
rect 513573 437868 513605 437902
rect 513639 437868 513674 437902
rect 513573 437812 513674 437868
rect 513573 437778 513605 437812
rect 513639 437778 513674 437812
rect 513573 437722 513674 437778
rect 513573 437688 513605 437722
rect 513639 437688 513674 437722
rect 513573 437632 513674 437688
rect 513573 437598 513605 437632
rect 513639 437598 513674 437632
rect 513573 437542 513674 437598
rect 513573 437508 513605 437542
rect 513639 437508 513674 437542
rect 513573 437452 513674 437508
rect 513573 437418 513605 437452
rect 513639 437418 513674 437452
rect 513573 437362 513674 437418
rect 512285 437295 512487 437328
rect 513573 437328 513605 437362
rect 513639 437328 513674 437362
rect 513573 437295 513674 437328
rect 503370 437261 513674 437295
rect 503370 437227 503486 437261
rect 503520 437227 503576 437261
rect 503610 437227 503666 437261
rect 503700 437227 503756 437261
rect 503790 437227 503846 437261
rect 503880 437227 503936 437261
rect 503970 437227 504026 437261
rect 504060 437227 504116 437261
rect 504150 437227 504206 437261
rect 504240 437227 504296 437261
rect 504330 437227 504386 437261
rect 504420 437227 504476 437261
rect 504510 437227 504566 437261
rect 504600 437227 504774 437261
rect 504808 437227 504864 437261
rect 504898 437227 504954 437261
rect 504988 437227 505044 437261
rect 505078 437227 505134 437261
rect 505168 437227 505224 437261
rect 505258 437227 505314 437261
rect 505348 437227 505404 437261
rect 505438 437227 505494 437261
rect 505528 437227 505584 437261
rect 505618 437227 505674 437261
rect 505708 437227 505764 437261
rect 505798 437227 505854 437261
rect 505888 437227 506062 437261
rect 506096 437227 506152 437261
rect 506186 437227 506242 437261
rect 506276 437227 506332 437261
rect 506366 437227 506422 437261
rect 506456 437227 506512 437261
rect 506546 437227 506602 437261
rect 506636 437227 506692 437261
rect 506726 437227 506782 437261
rect 506816 437227 506872 437261
rect 506906 437227 506962 437261
rect 506996 437227 507052 437261
rect 507086 437227 507142 437261
rect 507176 437227 507350 437261
rect 507384 437227 507440 437261
rect 507474 437227 507530 437261
rect 507564 437227 507620 437261
rect 507654 437227 507710 437261
rect 507744 437227 507800 437261
rect 507834 437227 507890 437261
rect 507924 437227 507980 437261
rect 508014 437227 508070 437261
rect 508104 437227 508160 437261
rect 508194 437227 508250 437261
rect 508284 437227 508340 437261
rect 508374 437227 508430 437261
rect 508464 437227 508638 437261
rect 508672 437227 508728 437261
rect 508762 437227 508818 437261
rect 508852 437227 508908 437261
rect 508942 437227 508998 437261
rect 509032 437227 509088 437261
rect 509122 437227 509178 437261
rect 509212 437227 509268 437261
rect 509302 437227 509358 437261
rect 509392 437227 509448 437261
rect 509482 437227 509538 437261
rect 509572 437227 509628 437261
rect 509662 437227 509718 437261
rect 509752 437227 509926 437261
rect 509960 437227 510016 437261
rect 510050 437227 510106 437261
rect 510140 437227 510196 437261
rect 510230 437227 510286 437261
rect 510320 437227 510376 437261
rect 510410 437227 510466 437261
rect 510500 437227 510556 437261
rect 510590 437227 510646 437261
rect 510680 437227 510736 437261
rect 510770 437227 510826 437261
rect 510860 437227 510916 437261
rect 510950 437227 511006 437261
rect 511040 437227 511214 437261
rect 511248 437227 511304 437261
rect 511338 437227 511394 437261
rect 511428 437227 511484 437261
rect 511518 437227 511574 437261
rect 511608 437227 511664 437261
rect 511698 437227 511754 437261
rect 511788 437227 511844 437261
rect 511878 437227 511934 437261
rect 511968 437227 512024 437261
rect 512058 437227 512114 437261
rect 512148 437227 512204 437261
rect 512238 437227 512294 437261
rect 512328 437227 512502 437261
rect 512536 437227 512592 437261
rect 512626 437227 512682 437261
rect 512716 437227 512772 437261
rect 512806 437227 512862 437261
rect 512896 437227 512952 437261
rect 512986 437227 513042 437261
rect 513076 437227 513132 437261
rect 513166 437227 513222 437261
rect 513256 437227 513312 437261
rect 513346 437227 513402 437261
rect 513436 437227 513492 437261
rect 513526 437227 513582 437261
rect 513616 437227 513674 437261
rect 503370 437160 513674 437227
rect 516598 437816 522950 437840
rect 516598 437246 516622 437816
rect 522926 437246 522950 437816
rect 516598 437222 522950 437246
rect 503370 437126 503486 437160
rect 503520 437126 503576 437160
rect 503610 437126 503666 437160
rect 503700 437126 503756 437160
rect 503790 437126 503846 437160
rect 503880 437126 503936 437160
rect 503970 437126 504026 437160
rect 504060 437126 504116 437160
rect 504150 437126 504206 437160
rect 504240 437126 504296 437160
rect 504330 437126 504386 437160
rect 504420 437126 504476 437160
rect 504510 437126 504566 437160
rect 504600 437126 504774 437160
rect 504808 437126 504864 437160
rect 504898 437126 504954 437160
rect 504988 437126 505044 437160
rect 505078 437126 505134 437160
rect 505168 437126 505224 437160
rect 505258 437126 505314 437160
rect 505348 437126 505404 437160
rect 505438 437126 505494 437160
rect 505528 437126 505584 437160
rect 505618 437126 505674 437160
rect 505708 437126 505764 437160
rect 505798 437126 505854 437160
rect 505888 437126 506062 437160
rect 506096 437126 506152 437160
rect 506186 437126 506242 437160
rect 506276 437126 506332 437160
rect 506366 437126 506422 437160
rect 506456 437126 506512 437160
rect 506546 437126 506602 437160
rect 506636 437126 506692 437160
rect 506726 437126 506782 437160
rect 506816 437126 506872 437160
rect 506906 437126 506962 437160
rect 506996 437126 507052 437160
rect 507086 437126 507142 437160
rect 507176 437126 507350 437160
rect 507384 437126 507440 437160
rect 507474 437126 507530 437160
rect 507564 437126 507620 437160
rect 507654 437126 507710 437160
rect 507744 437126 507800 437160
rect 507834 437126 507890 437160
rect 507924 437126 507980 437160
rect 508014 437126 508070 437160
rect 508104 437126 508160 437160
rect 508194 437126 508250 437160
rect 508284 437126 508340 437160
rect 508374 437126 508430 437160
rect 508464 437126 508638 437160
rect 508672 437126 508728 437160
rect 508762 437126 508818 437160
rect 508852 437126 508908 437160
rect 508942 437126 508998 437160
rect 509032 437126 509088 437160
rect 509122 437126 509178 437160
rect 509212 437126 509268 437160
rect 509302 437126 509358 437160
rect 509392 437126 509448 437160
rect 509482 437126 509538 437160
rect 509572 437126 509628 437160
rect 509662 437126 509718 437160
rect 509752 437126 509926 437160
rect 509960 437126 510016 437160
rect 510050 437126 510106 437160
rect 510140 437126 510196 437160
rect 510230 437126 510286 437160
rect 510320 437126 510376 437160
rect 510410 437126 510466 437160
rect 510500 437126 510556 437160
rect 510590 437126 510646 437160
rect 510680 437126 510736 437160
rect 510770 437126 510826 437160
rect 510860 437126 510916 437160
rect 510950 437126 511006 437160
rect 511040 437126 511214 437160
rect 511248 437126 511304 437160
rect 511338 437126 511394 437160
rect 511428 437126 511484 437160
rect 511518 437126 511574 437160
rect 511608 437126 511664 437160
rect 511698 437126 511754 437160
rect 511788 437126 511844 437160
rect 511878 437126 511934 437160
rect 511968 437126 512024 437160
rect 512058 437126 512114 437160
rect 512148 437126 512204 437160
rect 512238 437126 512294 437160
rect 512328 437126 512502 437160
rect 512536 437126 512592 437160
rect 512626 437126 512682 437160
rect 512716 437126 512772 437160
rect 512806 437126 512862 437160
rect 512896 437126 512952 437160
rect 512986 437126 513042 437160
rect 513076 437126 513132 437160
rect 513166 437126 513222 437160
rect 513256 437126 513312 437160
rect 513346 437126 513402 437160
rect 513436 437126 513492 437160
rect 513526 437126 513582 437160
rect 513616 437126 513674 437160
rect 503370 437093 513674 437126
rect 503370 437064 503471 437093
rect 503370 437030 503402 437064
rect 503436 437030 503471 437064
rect 504557 437064 504759 437093
rect 503370 436974 503471 437030
rect 503370 436940 503402 436974
rect 503436 436940 503471 436974
rect 503370 436884 503471 436940
rect 503370 436850 503402 436884
rect 503436 436850 503471 436884
rect 503370 436794 503471 436850
rect 503370 436760 503402 436794
rect 503436 436760 503471 436794
rect 503370 436704 503471 436760
rect 503370 436670 503402 436704
rect 503436 436670 503471 436704
rect 503370 436614 503471 436670
rect 503370 436580 503402 436614
rect 503436 436580 503471 436614
rect 503370 436524 503471 436580
rect 503370 436490 503402 436524
rect 503436 436490 503471 436524
rect 503370 436434 503471 436490
rect 503370 436400 503402 436434
rect 503436 436400 503471 436434
rect 503370 436344 503471 436400
rect 503370 436310 503402 436344
rect 503436 436310 503471 436344
rect 503370 436254 503471 436310
rect 503370 436220 503402 436254
rect 503436 436220 503471 436254
rect 503370 436164 503471 436220
rect 503370 436130 503402 436164
rect 503436 436130 503471 436164
rect 503370 436074 503471 436130
rect 503370 436040 503402 436074
rect 503436 436040 503471 436074
rect 504557 437030 504589 437064
rect 504623 437030 504690 437064
rect 504724 437030 504759 437064
rect 505845 437064 506047 437093
rect 504557 436974 504759 437030
rect 504557 436940 504589 436974
rect 504623 436940 504690 436974
rect 504724 436940 504759 436974
rect 504557 436884 504759 436940
rect 504557 436850 504589 436884
rect 504623 436850 504690 436884
rect 504724 436850 504759 436884
rect 504557 436794 504759 436850
rect 504557 436760 504589 436794
rect 504623 436760 504690 436794
rect 504724 436760 504759 436794
rect 504557 436704 504759 436760
rect 504557 436670 504589 436704
rect 504623 436670 504690 436704
rect 504724 436670 504759 436704
rect 504557 436614 504759 436670
rect 504557 436580 504589 436614
rect 504623 436580 504690 436614
rect 504724 436580 504759 436614
rect 504557 436524 504759 436580
rect 504557 436490 504589 436524
rect 504623 436490 504690 436524
rect 504724 436490 504759 436524
rect 504557 436434 504759 436490
rect 504557 436400 504589 436434
rect 504623 436400 504690 436434
rect 504724 436400 504759 436434
rect 504557 436344 504759 436400
rect 504557 436310 504589 436344
rect 504623 436310 504690 436344
rect 504724 436310 504759 436344
rect 504557 436254 504759 436310
rect 504557 436220 504589 436254
rect 504623 436220 504690 436254
rect 504724 436220 504759 436254
rect 504557 436164 504759 436220
rect 504557 436130 504589 436164
rect 504623 436130 504690 436164
rect 504724 436130 504759 436164
rect 504557 436074 504759 436130
rect 503370 436007 503471 436040
rect 504557 436040 504589 436074
rect 504623 436040 504690 436074
rect 504724 436040 504759 436074
rect 505845 437030 505877 437064
rect 505911 437030 505978 437064
rect 506012 437030 506047 437064
rect 507133 437064 507335 437093
rect 505845 436974 506047 437030
rect 505845 436940 505877 436974
rect 505911 436940 505978 436974
rect 506012 436940 506047 436974
rect 505845 436884 506047 436940
rect 505845 436850 505877 436884
rect 505911 436850 505978 436884
rect 506012 436850 506047 436884
rect 505845 436794 506047 436850
rect 505845 436760 505877 436794
rect 505911 436760 505978 436794
rect 506012 436760 506047 436794
rect 505845 436704 506047 436760
rect 505845 436670 505877 436704
rect 505911 436670 505978 436704
rect 506012 436670 506047 436704
rect 505845 436614 506047 436670
rect 505845 436580 505877 436614
rect 505911 436580 505978 436614
rect 506012 436580 506047 436614
rect 505845 436524 506047 436580
rect 505845 436490 505877 436524
rect 505911 436490 505978 436524
rect 506012 436490 506047 436524
rect 505845 436434 506047 436490
rect 505845 436400 505877 436434
rect 505911 436400 505978 436434
rect 506012 436400 506047 436434
rect 505845 436344 506047 436400
rect 505845 436310 505877 436344
rect 505911 436310 505978 436344
rect 506012 436310 506047 436344
rect 505845 436254 506047 436310
rect 505845 436220 505877 436254
rect 505911 436220 505978 436254
rect 506012 436220 506047 436254
rect 505845 436164 506047 436220
rect 505845 436130 505877 436164
rect 505911 436130 505978 436164
rect 506012 436130 506047 436164
rect 505845 436074 506047 436130
rect 504557 436007 504759 436040
rect 505845 436040 505877 436074
rect 505911 436040 505978 436074
rect 506012 436040 506047 436074
rect 507133 437030 507165 437064
rect 507199 437030 507266 437064
rect 507300 437030 507335 437064
rect 508421 437064 508623 437093
rect 507133 436974 507335 437030
rect 507133 436940 507165 436974
rect 507199 436940 507266 436974
rect 507300 436940 507335 436974
rect 507133 436884 507335 436940
rect 507133 436850 507165 436884
rect 507199 436850 507266 436884
rect 507300 436850 507335 436884
rect 507133 436794 507335 436850
rect 507133 436760 507165 436794
rect 507199 436760 507266 436794
rect 507300 436760 507335 436794
rect 507133 436704 507335 436760
rect 507133 436670 507165 436704
rect 507199 436670 507266 436704
rect 507300 436670 507335 436704
rect 507133 436614 507335 436670
rect 507133 436580 507165 436614
rect 507199 436580 507266 436614
rect 507300 436580 507335 436614
rect 507133 436524 507335 436580
rect 507133 436490 507165 436524
rect 507199 436490 507266 436524
rect 507300 436490 507335 436524
rect 507133 436434 507335 436490
rect 507133 436400 507165 436434
rect 507199 436400 507266 436434
rect 507300 436400 507335 436434
rect 507133 436344 507335 436400
rect 507133 436310 507165 436344
rect 507199 436310 507266 436344
rect 507300 436310 507335 436344
rect 507133 436254 507335 436310
rect 507133 436220 507165 436254
rect 507199 436220 507266 436254
rect 507300 436220 507335 436254
rect 507133 436164 507335 436220
rect 507133 436130 507165 436164
rect 507199 436130 507266 436164
rect 507300 436130 507335 436164
rect 507133 436074 507335 436130
rect 505845 436007 506047 436040
rect 507133 436040 507165 436074
rect 507199 436040 507266 436074
rect 507300 436040 507335 436074
rect 508421 437030 508453 437064
rect 508487 437030 508554 437064
rect 508588 437030 508623 437064
rect 509709 437064 509911 437093
rect 508421 436974 508623 437030
rect 508421 436940 508453 436974
rect 508487 436940 508554 436974
rect 508588 436940 508623 436974
rect 508421 436884 508623 436940
rect 508421 436850 508453 436884
rect 508487 436850 508554 436884
rect 508588 436850 508623 436884
rect 508421 436794 508623 436850
rect 508421 436760 508453 436794
rect 508487 436760 508554 436794
rect 508588 436760 508623 436794
rect 508421 436704 508623 436760
rect 508421 436670 508453 436704
rect 508487 436670 508554 436704
rect 508588 436670 508623 436704
rect 508421 436614 508623 436670
rect 508421 436580 508453 436614
rect 508487 436580 508554 436614
rect 508588 436580 508623 436614
rect 508421 436524 508623 436580
rect 508421 436490 508453 436524
rect 508487 436490 508554 436524
rect 508588 436490 508623 436524
rect 508421 436434 508623 436490
rect 508421 436400 508453 436434
rect 508487 436400 508554 436434
rect 508588 436400 508623 436434
rect 508421 436344 508623 436400
rect 508421 436310 508453 436344
rect 508487 436310 508554 436344
rect 508588 436310 508623 436344
rect 508421 436254 508623 436310
rect 508421 436220 508453 436254
rect 508487 436220 508554 436254
rect 508588 436220 508623 436254
rect 508421 436164 508623 436220
rect 508421 436130 508453 436164
rect 508487 436130 508554 436164
rect 508588 436130 508623 436164
rect 508421 436074 508623 436130
rect 507133 436007 507335 436040
rect 508421 436040 508453 436074
rect 508487 436040 508554 436074
rect 508588 436040 508623 436074
rect 509709 437030 509741 437064
rect 509775 437030 509842 437064
rect 509876 437030 509911 437064
rect 510997 437064 511199 437093
rect 509709 436974 509911 437030
rect 509709 436940 509741 436974
rect 509775 436940 509842 436974
rect 509876 436940 509911 436974
rect 509709 436884 509911 436940
rect 509709 436850 509741 436884
rect 509775 436850 509842 436884
rect 509876 436850 509911 436884
rect 509709 436794 509911 436850
rect 509709 436760 509741 436794
rect 509775 436760 509842 436794
rect 509876 436760 509911 436794
rect 509709 436704 509911 436760
rect 509709 436670 509741 436704
rect 509775 436670 509842 436704
rect 509876 436670 509911 436704
rect 509709 436614 509911 436670
rect 509709 436580 509741 436614
rect 509775 436580 509842 436614
rect 509876 436580 509911 436614
rect 509709 436524 509911 436580
rect 509709 436490 509741 436524
rect 509775 436490 509842 436524
rect 509876 436490 509911 436524
rect 509709 436434 509911 436490
rect 509709 436400 509741 436434
rect 509775 436400 509842 436434
rect 509876 436400 509911 436434
rect 509709 436344 509911 436400
rect 509709 436310 509741 436344
rect 509775 436310 509842 436344
rect 509876 436310 509911 436344
rect 509709 436254 509911 436310
rect 509709 436220 509741 436254
rect 509775 436220 509842 436254
rect 509876 436220 509911 436254
rect 509709 436164 509911 436220
rect 509709 436130 509741 436164
rect 509775 436130 509842 436164
rect 509876 436130 509911 436164
rect 509709 436074 509911 436130
rect 508421 436007 508623 436040
rect 509709 436040 509741 436074
rect 509775 436040 509842 436074
rect 509876 436040 509911 436074
rect 510997 437030 511029 437064
rect 511063 437030 511130 437064
rect 511164 437030 511199 437064
rect 512285 437064 512487 437093
rect 510997 436974 511199 437030
rect 510997 436940 511029 436974
rect 511063 436940 511130 436974
rect 511164 436940 511199 436974
rect 510997 436884 511199 436940
rect 510997 436850 511029 436884
rect 511063 436850 511130 436884
rect 511164 436850 511199 436884
rect 510997 436794 511199 436850
rect 510997 436760 511029 436794
rect 511063 436760 511130 436794
rect 511164 436760 511199 436794
rect 510997 436704 511199 436760
rect 510997 436670 511029 436704
rect 511063 436670 511130 436704
rect 511164 436670 511199 436704
rect 510997 436614 511199 436670
rect 510997 436580 511029 436614
rect 511063 436580 511130 436614
rect 511164 436580 511199 436614
rect 510997 436524 511199 436580
rect 510997 436490 511029 436524
rect 511063 436490 511130 436524
rect 511164 436490 511199 436524
rect 510997 436434 511199 436490
rect 510997 436400 511029 436434
rect 511063 436400 511130 436434
rect 511164 436400 511199 436434
rect 510997 436344 511199 436400
rect 510997 436310 511029 436344
rect 511063 436310 511130 436344
rect 511164 436310 511199 436344
rect 510997 436254 511199 436310
rect 510997 436220 511029 436254
rect 511063 436220 511130 436254
rect 511164 436220 511199 436254
rect 510997 436164 511199 436220
rect 510997 436130 511029 436164
rect 511063 436130 511130 436164
rect 511164 436130 511199 436164
rect 510997 436074 511199 436130
rect 509709 436007 509911 436040
rect 510997 436040 511029 436074
rect 511063 436040 511130 436074
rect 511164 436040 511199 436074
rect 512285 437030 512317 437064
rect 512351 437030 512418 437064
rect 512452 437030 512487 437064
rect 513573 437064 513674 437093
rect 512285 436974 512487 437030
rect 512285 436940 512317 436974
rect 512351 436940 512418 436974
rect 512452 436940 512487 436974
rect 512285 436884 512487 436940
rect 512285 436850 512317 436884
rect 512351 436850 512418 436884
rect 512452 436850 512487 436884
rect 512285 436794 512487 436850
rect 512285 436760 512317 436794
rect 512351 436760 512418 436794
rect 512452 436760 512487 436794
rect 512285 436704 512487 436760
rect 512285 436670 512317 436704
rect 512351 436670 512418 436704
rect 512452 436670 512487 436704
rect 512285 436614 512487 436670
rect 512285 436580 512317 436614
rect 512351 436580 512418 436614
rect 512452 436580 512487 436614
rect 512285 436524 512487 436580
rect 512285 436490 512317 436524
rect 512351 436490 512418 436524
rect 512452 436490 512487 436524
rect 512285 436434 512487 436490
rect 512285 436400 512317 436434
rect 512351 436400 512418 436434
rect 512452 436400 512487 436434
rect 512285 436344 512487 436400
rect 512285 436310 512317 436344
rect 512351 436310 512418 436344
rect 512452 436310 512487 436344
rect 512285 436254 512487 436310
rect 512285 436220 512317 436254
rect 512351 436220 512418 436254
rect 512452 436220 512487 436254
rect 512285 436164 512487 436220
rect 512285 436130 512317 436164
rect 512351 436130 512418 436164
rect 512452 436130 512487 436164
rect 512285 436074 512487 436130
rect 510997 436007 511199 436040
rect 512285 436040 512317 436074
rect 512351 436040 512418 436074
rect 512452 436040 512487 436074
rect 513573 437030 513605 437064
rect 513639 437030 513674 437064
rect 513573 436974 513674 437030
rect 513573 436940 513605 436974
rect 513639 436940 513674 436974
rect 513573 436884 513674 436940
rect 513573 436850 513605 436884
rect 513639 436850 513674 436884
rect 513573 436794 513674 436850
rect 513573 436760 513605 436794
rect 513639 436760 513674 436794
rect 513573 436704 513674 436760
rect 513573 436670 513605 436704
rect 513639 436670 513674 436704
rect 513573 436614 513674 436670
rect 513573 436580 513605 436614
rect 513639 436580 513674 436614
rect 513573 436524 513674 436580
rect 513573 436490 513605 436524
rect 513639 436490 513674 436524
rect 513573 436434 513674 436490
rect 513573 436400 513605 436434
rect 513639 436400 513674 436434
rect 513573 436344 513674 436400
rect 513573 436310 513605 436344
rect 513639 436310 513674 436344
rect 513573 436254 513674 436310
rect 513573 436220 513605 436254
rect 513639 436220 513674 436254
rect 513573 436164 513674 436220
rect 513573 436130 513605 436164
rect 513639 436130 513674 436164
rect 513573 436074 513674 436130
rect 512285 436007 512487 436040
rect 513573 436040 513605 436074
rect 513639 436040 513674 436074
rect 513573 436007 513674 436040
rect 503370 435973 513674 436007
rect 503370 435939 503486 435973
rect 503520 435939 503576 435973
rect 503610 435939 503666 435973
rect 503700 435939 503756 435973
rect 503790 435939 503846 435973
rect 503880 435939 503936 435973
rect 503970 435939 504026 435973
rect 504060 435939 504116 435973
rect 504150 435939 504206 435973
rect 504240 435939 504296 435973
rect 504330 435939 504386 435973
rect 504420 435939 504476 435973
rect 504510 435939 504566 435973
rect 504600 435939 504774 435973
rect 504808 435939 504864 435973
rect 504898 435939 504954 435973
rect 504988 435939 505044 435973
rect 505078 435939 505134 435973
rect 505168 435939 505224 435973
rect 505258 435939 505314 435973
rect 505348 435939 505404 435973
rect 505438 435939 505494 435973
rect 505528 435939 505584 435973
rect 505618 435939 505674 435973
rect 505708 435939 505764 435973
rect 505798 435939 505854 435973
rect 505888 435939 506062 435973
rect 506096 435939 506152 435973
rect 506186 435939 506242 435973
rect 506276 435939 506332 435973
rect 506366 435939 506422 435973
rect 506456 435939 506512 435973
rect 506546 435939 506602 435973
rect 506636 435939 506692 435973
rect 506726 435939 506782 435973
rect 506816 435939 506872 435973
rect 506906 435939 506962 435973
rect 506996 435939 507052 435973
rect 507086 435939 507142 435973
rect 507176 435939 507350 435973
rect 507384 435939 507440 435973
rect 507474 435939 507530 435973
rect 507564 435939 507620 435973
rect 507654 435939 507710 435973
rect 507744 435939 507800 435973
rect 507834 435939 507890 435973
rect 507924 435939 507980 435973
rect 508014 435939 508070 435973
rect 508104 435939 508160 435973
rect 508194 435939 508250 435973
rect 508284 435939 508340 435973
rect 508374 435939 508430 435973
rect 508464 435939 508638 435973
rect 508672 435939 508728 435973
rect 508762 435939 508818 435973
rect 508852 435939 508908 435973
rect 508942 435939 508998 435973
rect 509032 435939 509088 435973
rect 509122 435939 509178 435973
rect 509212 435939 509268 435973
rect 509302 435939 509358 435973
rect 509392 435939 509448 435973
rect 509482 435939 509538 435973
rect 509572 435939 509628 435973
rect 509662 435939 509718 435973
rect 509752 435939 509926 435973
rect 509960 435939 510016 435973
rect 510050 435939 510106 435973
rect 510140 435939 510196 435973
rect 510230 435939 510286 435973
rect 510320 435939 510376 435973
rect 510410 435939 510466 435973
rect 510500 435939 510556 435973
rect 510590 435939 510646 435973
rect 510680 435939 510736 435973
rect 510770 435939 510826 435973
rect 510860 435939 510916 435973
rect 510950 435939 511006 435973
rect 511040 435939 511214 435973
rect 511248 435939 511304 435973
rect 511338 435939 511394 435973
rect 511428 435939 511484 435973
rect 511518 435939 511574 435973
rect 511608 435939 511664 435973
rect 511698 435939 511754 435973
rect 511788 435939 511844 435973
rect 511878 435939 511934 435973
rect 511968 435939 512024 435973
rect 512058 435939 512114 435973
rect 512148 435939 512204 435973
rect 512238 435939 512294 435973
rect 512328 435939 512502 435973
rect 512536 435939 512592 435973
rect 512626 435939 512682 435973
rect 512716 435939 512772 435973
rect 512806 435939 512862 435973
rect 512896 435939 512952 435973
rect 512986 435939 513042 435973
rect 513076 435939 513132 435973
rect 513166 435939 513222 435973
rect 513256 435939 513312 435973
rect 513346 435939 513402 435973
rect 513436 435939 513492 435973
rect 513526 435939 513582 435973
rect 513616 435939 513674 435973
rect 503370 435872 513674 435939
rect 503370 435838 503486 435872
rect 503520 435838 503576 435872
rect 503610 435838 503666 435872
rect 503700 435838 503756 435872
rect 503790 435838 503846 435872
rect 503880 435838 503936 435872
rect 503970 435838 504026 435872
rect 504060 435838 504116 435872
rect 504150 435838 504206 435872
rect 504240 435838 504296 435872
rect 504330 435838 504386 435872
rect 504420 435838 504476 435872
rect 504510 435838 504566 435872
rect 504600 435838 504774 435872
rect 504808 435838 504864 435872
rect 504898 435838 504954 435872
rect 504988 435838 505044 435872
rect 505078 435838 505134 435872
rect 505168 435838 505224 435872
rect 505258 435838 505314 435872
rect 505348 435838 505404 435872
rect 505438 435838 505494 435872
rect 505528 435838 505584 435872
rect 505618 435838 505674 435872
rect 505708 435838 505764 435872
rect 505798 435838 505854 435872
rect 505888 435838 506062 435872
rect 506096 435838 506152 435872
rect 506186 435838 506242 435872
rect 506276 435838 506332 435872
rect 506366 435838 506422 435872
rect 506456 435838 506512 435872
rect 506546 435838 506602 435872
rect 506636 435838 506692 435872
rect 506726 435838 506782 435872
rect 506816 435838 506872 435872
rect 506906 435838 506962 435872
rect 506996 435838 507052 435872
rect 507086 435838 507142 435872
rect 507176 435838 507350 435872
rect 507384 435838 507440 435872
rect 507474 435838 507530 435872
rect 507564 435838 507620 435872
rect 507654 435838 507710 435872
rect 507744 435838 507800 435872
rect 507834 435838 507890 435872
rect 507924 435838 507980 435872
rect 508014 435838 508070 435872
rect 508104 435838 508160 435872
rect 508194 435838 508250 435872
rect 508284 435838 508340 435872
rect 508374 435838 508430 435872
rect 508464 435838 508638 435872
rect 508672 435838 508728 435872
rect 508762 435838 508818 435872
rect 508852 435838 508908 435872
rect 508942 435838 508998 435872
rect 509032 435838 509088 435872
rect 509122 435838 509178 435872
rect 509212 435838 509268 435872
rect 509302 435838 509358 435872
rect 509392 435838 509448 435872
rect 509482 435838 509538 435872
rect 509572 435838 509628 435872
rect 509662 435838 509718 435872
rect 509752 435838 509926 435872
rect 509960 435838 510016 435872
rect 510050 435838 510106 435872
rect 510140 435838 510196 435872
rect 510230 435838 510286 435872
rect 510320 435838 510376 435872
rect 510410 435838 510466 435872
rect 510500 435838 510556 435872
rect 510590 435838 510646 435872
rect 510680 435838 510736 435872
rect 510770 435838 510826 435872
rect 510860 435838 510916 435872
rect 510950 435838 511006 435872
rect 511040 435838 511214 435872
rect 511248 435838 511304 435872
rect 511338 435838 511394 435872
rect 511428 435838 511484 435872
rect 511518 435838 511574 435872
rect 511608 435838 511664 435872
rect 511698 435838 511754 435872
rect 511788 435838 511844 435872
rect 511878 435838 511934 435872
rect 511968 435838 512024 435872
rect 512058 435838 512114 435872
rect 512148 435838 512204 435872
rect 512238 435838 512294 435872
rect 512328 435838 512502 435872
rect 512536 435838 512592 435872
rect 512626 435838 512682 435872
rect 512716 435838 512772 435872
rect 512806 435838 512862 435872
rect 512896 435838 512952 435872
rect 512986 435838 513042 435872
rect 513076 435838 513132 435872
rect 513166 435838 513222 435872
rect 513256 435838 513312 435872
rect 513346 435838 513402 435872
rect 513436 435838 513492 435872
rect 513526 435838 513582 435872
rect 513616 435838 513674 435872
rect 503370 435805 513674 435838
rect 503370 435776 503471 435805
rect 503370 435742 503402 435776
rect 503436 435742 503471 435776
rect 504557 435776 504759 435805
rect 503370 435686 503471 435742
rect 503370 435652 503402 435686
rect 503436 435652 503471 435686
rect 503370 435596 503471 435652
rect 503370 435562 503402 435596
rect 503436 435562 503471 435596
rect 503370 435506 503471 435562
rect 503370 435472 503402 435506
rect 503436 435472 503471 435506
rect 503370 435416 503471 435472
rect 503370 435382 503402 435416
rect 503436 435382 503471 435416
rect 503370 435326 503471 435382
rect 503370 435292 503402 435326
rect 503436 435292 503471 435326
rect 503370 435236 503471 435292
rect 503370 435202 503402 435236
rect 503436 435202 503471 435236
rect 503370 435146 503471 435202
rect 503370 435112 503402 435146
rect 503436 435112 503471 435146
rect 503370 435056 503471 435112
rect 503370 435022 503402 435056
rect 503436 435022 503471 435056
rect 503370 434966 503471 435022
rect 503370 434932 503402 434966
rect 503436 434932 503471 434966
rect 503370 434876 503471 434932
rect 503370 434842 503402 434876
rect 503436 434842 503471 434876
rect 503370 434786 503471 434842
rect 503370 434752 503402 434786
rect 503436 434752 503471 434786
rect 504557 435742 504589 435776
rect 504623 435742 504690 435776
rect 504724 435742 504759 435776
rect 505845 435776 506047 435805
rect 504557 435686 504759 435742
rect 504557 435652 504589 435686
rect 504623 435652 504690 435686
rect 504724 435652 504759 435686
rect 504557 435596 504759 435652
rect 504557 435562 504589 435596
rect 504623 435562 504690 435596
rect 504724 435562 504759 435596
rect 504557 435506 504759 435562
rect 504557 435472 504589 435506
rect 504623 435472 504690 435506
rect 504724 435472 504759 435506
rect 504557 435416 504759 435472
rect 504557 435382 504589 435416
rect 504623 435382 504690 435416
rect 504724 435382 504759 435416
rect 504557 435326 504759 435382
rect 504557 435292 504589 435326
rect 504623 435292 504690 435326
rect 504724 435292 504759 435326
rect 504557 435236 504759 435292
rect 504557 435202 504589 435236
rect 504623 435202 504690 435236
rect 504724 435202 504759 435236
rect 504557 435146 504759 435202
rect 504557 435112 504589 435146
rect 504623 435112 504690 435146
rect 504724 435112 504759 435146
rect 504557 435056 504759 435112
rect 504557 435022 504589 435056
rect 504623 435022 504690 435056
rect 504724 435022 504759 435056
rect 504557 434966 504759 435022
rect 504557 434932 504589 434966
rect 504623 434932 504690 434966
rect 504724 434932 504759 434966
rect 504557 434876 504759 434932
rect 504557 434842 504589 434876
rect 504623 434842 504690 434876
rect 504724 434842 504759 434876
rect 504557 434786 504759 434842
rect 503370 434719 503471 434752
rect 504557 434752 504589 434786
rect 504623 434752 504690 434786
rect 504724 434752 504759 434786
rect 505845 435742 505877 435776
rect 505911 435742 505978 435776
rect 506012 435742 506047 435776
rect 507133 435776 507335 435805
rect 505845 435686 506047 435742
rect 505845 435652 505877 435686
rect 505911 435652 505978 435686
rect 506012 435652 506047 435686
rect 505845 435596 506047 435652
rect 505845 435562 505877 435596
rect 505911 435562 505978 435596
rect 506012 435562 506047 435596
rect 505845 435506 506047 435562
rect 505845 435472 505877 435506
rect 505911 435472 505978 435506
rect 506012 435472 506047 435506
rect 505845 435416 506047 435472
rect 505845 435382 505877 435416
rect 505911 435382 505978 435416
rect 506012 435382 506047 435416
rect 505845 435326 506047 435382
rect 505845 435292 505877 435326
rect 505911 435292 505978 435326
rect 506012 435292 506047 435326
rect 505845 435236 506047 435292
rect 505845 435202 505877 435236
rect 505911 435202 505978 435236
rect 506012 435202 506047 435236
rect 505845 435146 506047 435202
rect 505845 435112 505877 435146
rect 505911 435112 505978 435146
rect 506012 435112 506047 435146
rect 505845 435056 506047 435112
rect 505845 435022 505877 435056
rect 505911 435022 505978 435056
rect 506012 435022 506047 435056
rect 505845 434966 506047 435022
rect 505845 434932 505877 434966
rect 505911 434932 505978 434966
rect 506012 434932 506047 434966
rect 505845 434876 506047 434932
rect 505845 434842 505877 434876
rect 505911 434842 505978 434876
rect 506012 434842 506047 434876
rect 505845 434786 506047 434842
rect 504557 434719 504759 434752
rect 505845 434752 505877 434786
rect 505911 434752 505978 434786
rect 506012 434752 506047 434786
rect 507133 435742 507165 435776
rect 507199 435742 507266 435776
rect 507300 435742 507335 435776
rect 508421 435776 508623 435805
rect 507133 435686 507335 435742
rect 507133 435652 507165 435686
rect 507199 435652 507266 435686
rect 507300 435652 507335 435686
rect 507133 435596 507335 435652
rect 507133 435562 507165 435596
rect 507199 435562 507266 435596
rect 507300 435562 507335 435596
rect 507133 435506 507335 435562
rect 507133 435472 507165 435506
rect 507199 435472 507266 435506
rect 507300 435472 507335 435506
rect 507133 435416 507335 435472
rect 507133 435382 507165 435416
rect 507199 435382 507266 435416
rect 507300 435382 507335 435416
rect 507133 435326 507335 435382
rect 507133 435292 507165 435326
rect 507199 435292 507266 435326
rect 507300 435292 507335 435326
rect 507133 435236 507335 435292
rect 507133 435202 507165 435236
rect 507199 435202 507266 435236
rect 507300 435202 507335 435236
rect 507133 435146 507335 435202
rect 507133 435112 507165 435146
rect 507199 435112 507266 435146
rect 507300 435112 507335 435146
rect 507133 435056 507335 435112
rect 507133 435022 507165 435056
rect 507199 435022 507266 435056
rect 507300 435022 507335 435056
rect 507133 434966 507335 435022
rect 507133 434932 507165 434966
rect 507199 434932 507266 434966
rect 507300 434932 507335 434966
rect 507133 434876 507335 434932
rect 507133 434842 507165 434876
rect 507199 434842 507266 434876
rect 507300 434842 507335 434876
rect 507133 434786 507335 434842
rect 505845 434719 506047 434752
rect 507133 434752 507165 434786
rect 507199 434752 507266 434786
rect 507300 434752 507335 434786
rect 508421 435742 508453 435776
rect 508487 435742 508554 435776
rect 508588 435742 508623 435776
rect 509709 435776 509911 435805
rect 508421 435686 508623 435742
rect 508421 435652 508453 435686
rect 508487 435652 508554 435686
rect 508588 435652 508623 435686
rect 508421 435596 508623 435652
rect 508421 435562 508453 435596
rect 508487 435562 508554 435596
rect 508588 435562 508623 435596
rect 508421 435506 508623 435562
rect 508421 435472 508453 435506
rect 508487 435472 508554 435506
rect 508588 435472 508623 435506
rect 508421 435416 508623 435472
rect 508421 435382 508453 435416
rect 508487 435382 508554 435416
rect 508588 435382 508623 435416
rect 508421 435326 508623 435382
rect 508421 435292 508453 435326
rect 508487 435292 508554 435326
rect 508588 435292 508623 435326
rect 508421 435236 508623 435292
rect 508421 435202 508453 435236
rect 508487 435202 508554 435236
rect 508588 435202 508623 435236
rect 508421 435146 508623 435202
rect 508421 435112 508453 435146
rect 508487 435112 508554 435146
rect 508588 435112 508623 435146
rect 508421 435056 508623 435112
rect 508421 435022 508453 435056
rect 508487 435022 508554 435056
rect 508588 435022 508623 435056
rect 508421 434966 508623 435022
rect 508421 434932 508453 434966
rect 508487 434932 508554 434966
rect 508588 434932 508623 434966
rect 508421 434876 508623 434932
rect 508421 434842 508453 434876
rect 508487 434842 508554 434876
rect 508588 434842 508623 434876
rect 508421 434786 508623 434842
rect 507133 434719 507335 434752
rect 508421 434752 508453 434786
rect 508487 434752 508554 434786
rect 508588 434752 508623 434786
rect 509709 435742 509741 435776
rect 509775 435742 509842 435776
rect 509876 435742 509911 435776
rect 510997 435776 511199 435805
rect 509709 435686 509911 435742
rect 509709 435652 509741 435686
rect 509775 435652 509842 435686
rect 509876 435652 509911 435686
rect 509709 435596 509911 435652
rect 509709 435562 509741 435596
rect 509775 435562 509842 435596
rect 509876 435562 509911 435596
rect 509709 435506 509911 435562
rect 509709 435472 509741 435506
rect 509775 435472 509842 435506
rect 509876 435472 509911 435506
rect 509709 435416 509911 435472
rect 509709 435382 509741 435416
rect 509775 435382 509842 435416
rect 509876 435382 509911 435416
rect 509709 435326 509911 435382
rect 509709 435292 509741 435326
rect 509775 435292 509842 435326
rect 509876 435292 509911 435326
rect 509709 435236 509911 435292
rect 509709 435202 509741 435236
rect 509775 435202 509842 435236
rect 509876 435202 509911 435236
rect 509709 435146 509911 435202
rect 509709 435112 509741 435146
rect 509775 435112 509842 435146
rect 509876 435112 509911 435146
rect 509709 435056 509911 435112
rect 509709 435022 509741 435056
rect 509775 435022 509842 435056
rect 509876 435022 509911 435056
rect 509709 434966 509911 435022
rect 509709 434932 509741 434966
rect 509775 434932 509842 434966
rect 509876 434932 509911 434966
rect 509709 434876 509911 434932
rect 509709 434842 509741 434876
rect 509775 434842 509842 434876
rect 509876 434842 509911 434876
rect 509709 434786 509911 434842
rect 508421 434719 508623 434752
rect 509709 434752 509741 434786
rect 509775 434752 509842 434786
rect 509876 434752 509911 434786
rect 510997 435742 511029 435776
rect 511063 435742 511130 435776
rect 511164 435742 511199 435776
rect 512285 435776 512487 435805
rect 510997 435686 511199 435742
rect 510997 435652 511029 435686
rect 511063 435652 511130 435686
rect 511164 435652 511199 435686
rect 510997 435596 511199 435652
rect 510997 435562 511029 435596
rect 511063 435562 511130 435596
rect 511164 435562 511199 435596
rect 510997 435506 511199 435562
rect 510997 435472 511029 435506
rect 511063 435472 511130 435506
rect 511164 435472 511199 435506
rect 510997 435416 511199 435472
rect 510997 435382 511029 435416
rect 511063 435382 511130 435416
rect 511164 435382 511199 435416
rect 510997 435326 511199 435382
rect 510997 435292 511029 435326
rect 511063 435292 511130 435326
rect 511164 435292 511199 435326
rect 510997 435236 511199 435292
rect 510997 435202 511029 435236
rect 511063 435202 511130 435236
rect 511164 435202 511199 435236
rect 510997 435146 511199 435202
rect 510997 435112 511029 435146
rect 511063 435112 511130 435146
rect 511164 435112 511199 435146
rect 510997 435056 511199 435112
rect 510997 435022 511029 435056
rect 511063 435022 511130 435056
rect 511164 435022 511199 435056
rect 510997 434966 511199 435022
rect 510997 434932 511029 434966
rect 511063 434932 511130 434966
rect 511164 434932 511199 434966
rect 510997 434876 511199 434932
rect 510997 434842 511029 434876
rect 511063 434842 511130 434876
rect 511164 434842 511199 434876
rect 510997 434786 511199 434842
rect 509709 434719 509911 434752
rect 510997 434752 511029 434786
rect 511063 434752 511130 434786
rect 511164 434752 511199 434786
rect 512285 435742 512317 435776
rect 512351 435742 512418 435776
rect 512452 435742 512487 435776
rect 513573 435776 513674 435805
rect 512285 435686 512487 435742
rect 512285 435652 512317 435686
rect 512351 435652 512418 435686
rect 512452 435652 512487 435686
rect 512285 435596 512487 435652
rect 512285 435562 512317 435596
rect 512351 435562 512418 435596
rect 512452 435562 512487 435596
rect 512285 435506 512487 435562
rect 512285 435472 512317 435506
rect 512351 435472 512418 435506
rect 512452 435472 512487 435506
rect 512285 435416 512487 435472
rect 512285 435382 512317 435416
rect 512351 435382 512418 435416
rect 512452 435382 512487 435416
rect 512285 435326 512487 435382
rect 512285 435292 512317 435326
rect 512351 435292 512418 435326
rect 512452 435292 512487 435326
rect 512285 435236 512487 435292
rect 512285 435202 512317 435236
rect 512351 435202 512418 435236
rect 512452 435202 512487 435236
rect 512285 435146 512487 435202
rect 512285 435112 512317 435146
rect 512351 435112 512418 435146
rect 512452 435112 512487 435146
rect 512285 435056 512487 435112
rect 512285 435022 512317 435056
rect 512351 435022 512418 435056
rect 512452 435022 512487 435056
rect 512285 434966 512487 435022
rect 512285 434932 512317 434966
rect 512351 434932 512418 434966
rect 512452 434932 512487 434966
rect 512285 434876 512487 434932
rect 512285 434842 512317 434876
rect 512351 434842 512418 434876
rect 512452 434842 512487 434876
rect 512285 434786 512487 434842
rect 510997 434719 511199 434752
rect 512285 434752 512317 434786
rect 512351 434752 512418 434786
rect 512452 434752 512487 434786
rect 513573 435742 513605 435776
rect 513639 435742 513674 435776
rect 513573 435686 513674 435742
rect 513573 435652 513605 435686
rect 513639 435652 513674 435686
rect 513573 435596 513674 435652
rect 513573 435562 513605 435596
rect 513639 435562 513674 435596
rect 513573 435506 513674 435562
rect 513573 435472 513605 435506
rect 513639 435472 513674 435506
rect 513573 435416 513674 435472
rect 513573 435382 513605 435416
rect 513639 435382 513674 435416
rect 513573 435326 513674 435382
rect 513573 435292 513605 435326
rect 513639 435292 513674 435326
rect 513573 435236 513674 435292
rect 513573 435202 513605 435236
rect 513639 435202 513674 435236
rect 513573 435146 513674 435202
rect 513573 435112 513605 435146
rect 513639 435112 513674 435146
rect 513573 435056 513674 435112
rect 513573 435022 513605 435056
rect 513639 435022 513674 435056
rect 513573 434966 513674 435022
rect 513573 434932 513605 434966
rect 513639 434932 513674 434966
rect 513573 434876 513674 434932
rect 513573 434842 513605 434876
rect 513639 434842 513674 434876
rect 513573 434786 513674 434842
rect 512285 434719 512487 434752
rect 513573 434752 513605 434786
rect 513639 434752 513674 434786
rect 513573 434719 513674 434752
rect 503370 434685 513674 434719
rect 503370 434651 503486 434685
rect 503520 434651 503576 434685
rect 503610 434651 503666 434685
rect 503700 434651 503756 434685
rect 503790 434651 503846 434685
rect 503880 434651 503936 434685
rect 503970 434651 504026 434685
rect 504060 434651 504116 434685
rect 504150 434651 504206 434685
rect 504240 434651 504296 434685
rect 504330 434651 504386 434685
rect 504420 434651 504476 434685
rect 504510 434651 504566 434685
rect 504600 434651 504774 434685
rect 504808 434651 504864 434685
rect 504898 434651 504954 434685
rect 504988 434651 505044 434685
rect 505078 434651 505134 434685
rect 505168 434651 505224 434685
rect 505258 434651 505314 434685
rect 505348 434651 505404 434685
rect 505438 434651 505494 434685
rect 505528 434651 505584 434685
rect 505618 434651 505674 434685
rect 505708 434651 505764 434685
rect 505798 434651 505854 434685
rect 505888 434651 506062 434685
rect 506096 434651 506152 434685
rect 506186 434651 506242 434685
rect 506276 434651 506332 434685
rect 506366 434651 506422 434685
rect 506456 434651 506512 434685
rect 506546 434651 506602 434685
rect 506636 434651 506692 434685
rect 506726 434651 506782 434685
rect 506816 434651 506872 434685
rect 506906 434651 506962 434685
rect 506996 434651 507052 434685
rect 507086 434651 507142 434685
rect 507176 434651 507350 434685
rect 507384 434651 507440 434685
rect 507474 434651 507530 434685
rect 507564 434651 507620 434685
rect 507654 434651 507710 434685
rect 507744 434651 507800 434685
rect 507834 434651 507890 434685
rect 507924 434651 507980 434685
rect 508014 434651 508070 434685
rect 508104 434651 508160 434685
rect 508194 434651 508250 434685
rect 508284 434651 508340 434685
rect 508374 434651 508430 434685
rect 508464 434651 508638 434685
rect 508672 434651 508728 434685
rect 508762 434651 508818 434685
rect 508852 434651 508908 434685
rect 508942 434651 508998 434685
rect 509032 434651 509088 434685
rect 509122 434651 509178 434685
rect 509212 434651 509268 434685
rect 509302 434651 509358 434685
rect 509392 434651 509448 434685
rect 509482 434651 509538 434685
rect 509572 434651 509628 434685
rect 509662 434651 509718 434685
rect 509752 434651 509926 434685
rect 509960 434651 510016 434685
rect 510050 434651 510106 434685
rect 510140 434651 510196 434685
rect 510230 434651 510286 434685
rect 510320 434651 510376 434685
rect 510410 434651 510466 434685
rect 510500 434651 510556 434685
rect 510590 434651 510646 434685
rect 510680 434651 510736 434685
rect 510770 434651 510826 434685
rect 510860 434651 510916 434685
rect 510950 434651 511006 434685
rect 511040 434651 511214 434685
rect 511248 434651 511304 434685
rect 511338 434651 511394 434685
rect 511428 434651 511484 434685
rect 511518 434651 511574 434685
rect 511608 434651 511664 434685
rect 511698 434651 511754 434685
rect 511788 434651 511844 434685
rect 511878 434651 511934 434685
rect 511968 434651 512024 434685
rect 512058 434651 512114 434685
rect 512148 434651 512204 434685
rect 512238 434651 512294 434685
rect 512328 434651 512502 434685
rect 512536 434651 512592 434685
rect 512626 434651 512682 434685
rect 512716 434651 512772 434685
rect 512806 434651 512862 434685
rect 512896 434651 512952 434685
rect 512986 434651 513042 434685
rect 513076 434651 513132 434685
rect 513166 434651 513222 434685
rect 513256 434651 513312 434685
rect 513346 434651 513402 434685
rect 513436 434651 513492 434685
rect 513526 434651 513582 434685
rect 513616 434651 513674 434685
rect 503370 434584 513674 434651
rect 503370 434550 503486 434584
rect 503520 434550 503576 434584
rect 503610 434550 503666 434584
rect 503700 434550 503756 434584
rect 503790 434550 503846 434584
rect 503880 434550 503936 434584
rect 503970 434550 504026 434584
rect 504060 434550 504116 434584
rect 504150 434550 504206 434584
rect 504240 434550 504296 434584
rect 504330 434550 504386 434584
rect 504420 434550 504476 434584
rect 504510 434550 504566 434584
rect 504600 434550 504774 434584
rect 504808 434550 504864 434584
rect 504898 434550 504954 434584
rect 504988 434550 505044 434584
rect 505078 434550 505134 434584
rect 505168 434550 505224 434584
rect 505258 434550 505314 434584
rect 505348 434550 505404 434584
rect 505438 434550 505494 434584
rect 505528 434550 505584 434584
rect 505618 434550 505674 434584
rect 505708 434550 505764 434584
rect 505798 434550 505854 434584
rect 505888 434550 506062 434584
rect 506096 434550 506152 434584
rect 506186 434550 506242 434584
rect 506276 434550 506332 434584
rect 506366 434550 506422 434584
rect 506456 434550 506512 434584
rect 506546 434550 506602 434584
rect 506636 434550 506692 434584
rect 506726 434550 506782 434584
rect 506816 434550 506872 434584
rect 506906 434550 506962 434584
rect 506996 434550 507052 434584
rect 507086 434550 507142 434584
rect 507176 434550 507350 434584
rect 507384 434550 507440 434584
rect 507474 434550 507530 434584
rect 507564 434550 507620 434584
rect 507654 434550 507710 434584
rect 507744 434550 507800 434584
rect 507834 434550 507890 434584
rect 507924 434550 507980 434584
rect 508014 434550 508070 434584
rect 508104 434550 508160 434584
rect 508194 434550 508250 434584
rect 508284 434550 508340 434584
rect 508374 434550 508430 434584
rect 508464 434550 508638 434584
rect 508672 434550 508728 434584
rect 508762 434550 508818 434584
rect 508852 434550 508908 434584
rect 508942 434550 508998 434584
rect 509032 434550 509088 434584
rect 509122 434550 509178 434584
rect 509212 434550 509268 434584
rect 509302 434550 509358 434584
rect 509392 434550 509448 434584
rect 509482 434550 509538 434584
rect 509572 434550 509628 434584
rect 509662 434550 509718 434584
rect 509752 434550 509926 434584
rect 509960 434550 510016 434584
rect 510050 434550 510106 434584
rect 510140 434550 510196 434584
rect 510230 434550 510286 434584
rect 510320 434550 510376 434584
rect 510410 434550 510466 434584
rect 510500 434550 510556 434584
rect 510590 434550 510646 434584
rect 510680 434550 510736 434584
rect 510770 434550 510826 434584
rect 510860 434550 510916 434584
rect 510950 434550 511006 434584
rect 511040 434550 511214 434584
rect 511248 434550 511304 434584
rect 511338 434550 511394 434584
rect 511428 434550 511484 434584
rect 511518 434550 511574 434584
rect 511608 434550 511664 434584
rect 511698 434550 511754 434584
rect 511788 434550 511844 434584
rect 511878 434550 511934 434584
rect 511968 434550 512024 434584
rect 512058 434550 512114 434584
rect 512148 434550 512204 434584
rect 512238 434550 512294 434584
rect 512328 434550 512502 434584
rect 512536 434550 512592 434584
rect 512626 434550 512682 434584
rect 512716 434550 512772 434584
rect 512806 434550 512862 434584
rect 512896 434550 512952 434584
rect 512986 434550 513042 434584
rect 513076 434550 513132 434584
rect 513166 434550 513222 434584
rect 513256 434550 513312 434584
rect 513346 434550 513402 434584
rect 513436 434550 513492 434584
rect 513526 434550 513582 434584
rect 513616 434550 513674 434584
rect 503370 434517 513674 434550
rect 503370 434488 503471 434517
rect 503370 434454 503402 434488
rect 503436 434454 503471 434488
rect 504557 434488 504759 434517
rect 503370 434398 503471 434454
rect 503370 434364 503402 434398
rect 503436 434364 503471 434398
rect 503370 434308 503471 434364
rect 503370 434274 503402 434308
rect 503436 434274 503471 434308
rect 503370 434218 503471 434274
rect 503370 434184 503402 434218
rect 503436 434184 503471 434218
rect 503370 434128 503471 434184
rect 503370 434094 503402 434128
rect 503436 434094 503471 434128
rect 503370 434038 503471 434094
rect 503370 434004 503402 434038
rect 503436 434004 503471 434038
rect 503370 433948 503471 434004
rect 503370 433914 503402 433948
rect 503436 433914 503471 433948
rect 503370 433858 503471 433914
rect 503370 433824 503402 433858
rect 503436 433824 503471 433858
rect 503370 433768 503471 433824
rect 503370 433734 503402 433768
rect 503436 433734 503471 433768
rect 503370 433678 503471 433734
rect 503370 433644 503402 433678
rect 503436 433644 503471 433678
rect 503370 433588 503471 433644
rect 503370 433554 503402 433588
rect 503436 433554 503471 433588
rect 503370 433498 503471 433554
rect 503370 433464 503402 433498
rect 503436 433464 503471 433498
rect 504557 434454 504589 434488
rect 504623 434454 504690 434488
rect 504724 434454 504759 434488
rect 505845 434488 506047 434517
rect 504557 434398 504759 434454
rect 504557 434364 504589 434398
rect 504623 434364 504690 434398
rect 504724 434364 504759 434398
rect 504557 434308 504759 434364
rect 504557 434274 504589 434308
rect 504623 434274 504690 434308
rect 504724 434274 504759 434308
rect 504557 434218 504759 434274
rect 504557 434184 504589 434218
rect 504623 434184 504690 434218
rect 504724 434184 504759 434218
rect 504557 434128 504759 434184
rect 504557 434094 504589 434128
rect 504623 434094 504690 434128
rect 504724 434094 504759 434128
rect 504557 434038 504759 434094
rect 504557 434004 504589 434038
rect 504623 434004 504690 434038
rect 504724 434004 504759 434038
rect 504557 433948 504759 434004
rect 504557 433914 504589 433948
rect 504623 433914 504690 433948
rect 504724 433914 504759 433948
rect 504557 433858 504759 433914
rect 504557 433824 504589 433858
rect 504623 433824 504690 433858
rect 504724 433824 504759 433858
rect 504557 433768 504759 433824
rect 504557 433734 504589 433768
rect 504623 433734 504690 433768
rect 504724 433734 504759 433768
rect 504557 433678 504759 433734
rect 504557 433644 504589 433678
rect 504623 433644 504690 433678
rect 504724 433644 504759 433678
rect 504557 433588 504759 433644
rect 504557 433554 504589 433588
rect 504623 433554 504690 433588
rect 504724 433554 504759 433588
rect 504557 433498 504759 433554
rect 503370 433431 503471 433464
rect 504557 433464 504589 433498
rect 504623 433464 504690 433498
rect 504724 433464 504759 433498
rect 505845 434454 505877 434488
rect 505911 434454 505978 434488
rect 506012 434454 506047 434488
rect 507133 434488 507335 434517
rect 505845 434398 506047 434454
rect 505845 434364 505877 434398
rect 505911 434364 505978 434398
rect 506012 434364 506047 434398
rect 505845 434308 506047 434364
rect 505845 434274 505877 434308
rect 505911 434274 505978 434308
rect 506012 434274 506047 434308
rect 505845 434218 506047 434274
rect 505845 434184 505877 434218
rect 505911 434184 505978 434218
rect 506012 434184 506047 434218
rect 505845 434128 506047 434184
rect 505845 434094 505877 434128
rect 505911 434094 505978 434128
rect 506012 434094 506047 434128
rect 505845 434038 506047 434094
rect 505845 434004 505877 434038
rect 505911 434004 505978 434038
rect 506012 434004 506047 434038
rect 505845 433948 506047 434004
rect 505845 433914 505877 433948
rect 505911 433914 505978 433948
rect 506012 433914 506047 433948
rect 505845 433858 506047 433914
rect 505845 433824 505877 433858
rect 505911 433824 505978 433858
rect 506012 433824 506047 433858
rect 505845 433768 506047 433824
rect 505845 433734 505877 433768
rect 505911 433734 505978 433768
rect 506012 433734 506047 433768
rect 505845 433678 506047 433734
rect 505845 433644 505877 433678
rect 505911 433644 505978 433678
rect 506012 433644 506047 433678
rect 505845 433588 506047 433644
rect 505845 433554 505877 433588
rect 505911 433554 505978 433588
rect 506012 433554 506047 433588
rect 505845 433498 506047 433554
rect 504557 433431 504759 433464
rect 505845 433464 505877 433498
rect 505911 433464 505978 433498
rect 506012 433464 506047 433498
rect 507133 434454 507165 434488
rect 507199 434454 507266 434488
rect 507300 434454 507335 434488
rect 508421 434488 508623 434517
rect 507133 434398 507335 434454
rect 507133 434364 507165 434398
rect 507199 434364 507266 434398
rect 507300 434364 507335 434398
rect 507133 434308 507335 434364
rect 507133 434274 507165 434308
rect 507199 434274 507266 434308
rect 507300 434274 507335 434308
rect 507133 434218 507335 434274
rect 507133 434184 507165 434218
rect 507199 434184 507266 434218
rect 507300 434184 507335 434218
rect 507133 434128 507335 434184
rect 507133 434094 507165 434128
rect 507199 434094 507266 434128
rect 507300 434094 507335 434128
rect 507133 434038 507335 434094
rect 507133 434004 507165 434038
rect 507199 434004 507266 434038
rect 507300 434004 507335 434038
rect 507133 433948 507335 434004
rect 507133 433914 507165 433948
rect 507199 433914 507266 433948
rect 507300 433914 507335 433948
rect 507133 433858 507335 433914
rect 507133 433824 507165 433858
rect 507199 433824 507266 433858
rect 507300 433824 507335 433858
rect 507133 433768 507335 433824
rect 507133 433734 507165 433768
rect 507199 433734 507266 433768
rect 507300 433734 507335 433768
rect 507133 433678 507335 433734
rect 507133 433644 507165 433678
rect 507199 433644 507266 433678
rect 507300 433644 507335 433678
rect 507133 433588 507335 433644
rect 507133 433554 507165 433588
rect 507199 433554 507266 433588
rect 507300 433554 507335 433588
rect 507133 433498 507335 433554
rect 505845 433431 506047 433464
rect 507133 433464 507165 433498
rect 507199 433464 507266 433498
rect 507300 433464 507335 433498
rect 508421 434454 508453 434488
rect 508487 434454 508554 434488
rect 508588 434454 508623 434488
rect 509709 434488 509911 434517
rect 508421 434398 508623 434454
rect 508421 434364 508453 434398
rect 508487 434364 508554 434398
rect 508588 434364 508623 434398
rect 508421 434308 508623 434364
rect 508421 434274 508453 434308
rect 508487 434274 508554 434308
rect 508588 434274 508623 434308
rect 508421 434218 508623 434274
rect 508421 434184 508453 434218
rect 508487 434184 508554 434218
rect 508588 434184 508623 434218
rect 508421 434128 508623 434184
rect 508421 434094 508453 434128
rect 508487 434094 508554 434128
rect 508588 434094 508623 434128
rect 508421 434038 508623 434094
rect 508421 434004 508453 434038
rect 508487 434004 508554 434038
rect 508588 434004 508623 434038
rect 508421 433948 508623 434004
rect 508421 433914 508453 433948
rect 508487 433914 508554 433948
rect 508588 433914 508623 433948
rect 508421 433858 508623 433914
rect 508421 433824 508453 433858
rect 508487 433824 508554 433858
rect 508588 433824 508623 433858
rect 508421 433768 508623 433824
rect 508421 433734 508453 433768
rect 508487 433734 508554 433768
rect 508588 433734 508623 433768
rect 508421 433678 508623 433734
rect 508421 433644 508453 433678
rect 508487 433644 508554 433678
rect 508588 433644 508623 433678
rect 508421 433588 508623 433644
rect 508421 433554 508453 433588
rect 508487 433554 508554 433588
rect 508588 433554 508623 433588
rect 508421 433498 508623 433554
rect 507133 433431 507335 433464
rect 508421 433464 508453 433498
rect 508487 433464 508554 433498
rect 508588 433464 508623 433498
rect 509709 434454 509741 434488
rect 509775 434454 509842 434488
rect 509876 434454 509911 434488
rect 510997 434488 511199 434517
rect 509709 434398 509911 434454
rect 509709 434364 509741 434398
rect 509775 434364 509842 434398
rect 509876 434364 509911 434398
rect 509709 434308 509911 434364
rect 509709 434274 509741 434308
rect 509775 434274 509842 434308
rect 509876 434274 509911 434308
rect 509709 434218 509911 434274
rect 509709 434184 509741 434218
rect 509775 434184 509842 434218
rect 509876 434184 509911 434218
rect 509709 434128 509911 434184
rect 509709 434094 509741 434128
rect 509775 434094 509842 434128
rect 509876 434094 509911 434128
rect 509709 434038 509911 434094
rect 509709 434004 509741 434038
rect 509775 434004 509842 434038
rect 509876 434004 509911 434038
rect 509709 433948 509911 434004
rect 509709 433914 509741 433948
rect 509775 433914 509842 433948
rect 509876 433914 509911 433948
rect 509709 433858 509911 433914
rect 509709 433824 509741 433858
rect 509775 433824 509842 433858
rect 509876 433824 509911 433858
rect 509709 433768 509911 433824
rect 509709 433734 509741 433768
rect 509775 433734 509842 433768
rect 509876 433734 509911 433768
rect 509709 433678 509911 433734
rect 509709 433644 509741 433678
rect 509775 433644 509842 433678
rect 509876 433644 509911 433678
rect 509709 433588 509911 433644
rect 509709 433554 509741 433588
rect 509775 433554 509842 433588
rect 509876 433554 509911 433588
rect 509709 433498 509911 433554
rect 508421 433431 508623 433464
rect 509709 433464 509741 433498
rect 509775 433464 509842 433498
rect 509876 433464 509911 433498
rect 510997 434454 511029 434488
rect 511063 434454 511130 434488
rect 511164 434454 511199 434488
rect 512285 434488 512487 434517
rect 510997 434398 511199 434454
rect 510997 434364 511029 434398
rect 511063 434364 511130 434398
rect 511164 434364 511199 434398
rect 510997 434308 511199 434364
rect 510997 434274 511029 434308
rect 511063 434274 511130 434308
rect 511164 434274 511199 434308
rect 510997 434218 511199 434274
rect 510997 434184 511029 434218
rect 511063 434184 511130 434218
rect 511164 434184 511199 434218
rect 510997 434128 511199 434184
rect 510997 434094 511029 434128
rect 511063 434094 511130 434128
rect 511164 434094 511199 434128
rect 510997 434038 511199 434094
rect 510997 434004 511029 434038
rect 511063 434004 511130 434038
rect 511164 434004 511199 434038
rect 510997 433948 511199 434004
rect 510997 433914 511029 433948
rect 511063 433914 511130 433948
rect 511164 433914 511199 433948
rect 510997 433858 511199 433914
rect 510997 433824 511029 433858
rect 511063 433824 511130 433858
rect 511164 433824 511199 433858
rect 510997 433768 511199 433824
rect 510997 433734 511029 433768
rect 511063 433734 511130 433768
rect 511164 433734 511199 433768
rect 510997 433678 511199 433734
rect 510997 433644 511029 433678
rect 511063 433644 511130 433678
rect 511164 433644 511199 433678
rect 510997 433588 511199 433644
rect 510997 433554 511029 433588
rect 511063 433554 511130 433588
rect 511164 433554 511199 433588
rect 510997 433498 511199 433554
rect 509709 433431 509911 433464
rect 510997 433464 511029 433498
rect 511063 433464 511130 433498
rect 511164 433464 511199 433498
rect 512285 434454 512317 434488
rect 512351 434454 512418 434488
rect 512452 434454 512487 434488
rect 513573 434488 513674 434517
rect 512285 434398 512487 434454
rect 512285 434364 512317 434398
rect 512351 434364 512418 434398
rect 512452 434364 512487 434398
rect 512285 434308 512487 434364
rect 512285 434274 512317 434308
rect 512351 434274 512418 434308
rect 512452 434274 512487 434308
rect 512285 434218 512487 434274
rect 512285 434184 512317 434218
rect 512351 434184 512418 434218
rect 512452 434184 512487 434218
rect 512285 434128 512487 434184
rect 512285 434094 512317 434128
rect 512351 434094 512418 434128
rect 512452 434094 512487 434128
rect 512285 434038 512487 434094
rect 512285 434004 512317 434038
rect 512351 434004 512418 434038
rect 512452 434004 512487 434038
rect 512285 433948 512487 434004
rect 512285 433914 512317 433948
rect 512351 433914 512418 433948
rect 512452 433914 512487 433948
rect 512285 433858 512487 433914
rect 512285 433824 512317 433858
rect 512351 433824 512418 433858
rect 512452 433824 512487 433858
rect 512285 433768 512487 433824
rect 512285 433734 512317 433768
rect 512351 433734 512418 433768
rect 512452 433734 512487 433768
rect 512285 433678 512487 433734
rect 512285 433644 512317 433678
rect 512351 433644 512418 433678
rect 512452 433644 512487 433678
rect 512285 433588 512487 433644
rect 512285 433554 512317 433588
rect 512351 433554 512418 433588
rect 512452 433554 512487 433588
rect 512285 433498 512487 433554
rect 510997 433431 511199 433464
rect 512285 433464 512317 433498
rect 512351 433464 512418 433498
rect 512452 433464 512487 433498
rect 513573 434454 513605 434488
rect 513639 434454 513674 434488
rect 513573 434398 513674 434454
rect 513573 434364 513605 434398
rect 513639 434364 513674 434398
rect 513573 434308 513674 434364
rect 513573 434274 513605 434308
rect 513639 434274 513674 434308
rect 513573 434218 513674 434274
rect 513573 434184 513605 434218
rect 513639 434184 513674 434218
rect 513573 434128 513674 434184
rect 513573 434094 513605 434128
rect 513639 434094 513674 434128
rect 513573 434038 513674 434094
rect 513573 434004 513605 434038
rect 513639 434004 513674 434038
rect 513573 433948 513674 434004
rect 513573 433914 513605 433948
rect 513639 433914 513674 433948
rect 513573 433858 513674 433914
rect 513573 433824 513605 433858
rect 513639 433824 513674 433858
rect 513573 433768 513674 433824
rect 513573 433734 513605 433768
rect 513639 433734 513674 433768
rect 513573 433678 513674 433734
rect 513573 433644 513605 433678
rect 513639 433644 513674 433678
rect 513573 433588 513674 433644
rect 513573 433554 513605 433588
rect 513639 433554 513674 433588
rect 513573 433498 513674 433554
rect 512285 433431 512487 433464
rect 513573 433464 513605 433498
rect 513639 433464 513674 433498
rect 513573 433431 513674 433464
rect 503370 433397 513674 433431
rect 503370 433363 503486 433397
rect 503520 433363 503576 433397
rect 503610 433363 503666 433397
rect 503700 433363 503756 433397
rect 503790 433363 503846 433397
rect 503880 433363 503936 433397
rect 503970 433363 504026 433397
rect 504060 433363 504116 433397
rect 504150 433363 504206 433397
rect 504240 433363 504296 433397
rect 504330 433363 504386 433397
rect 504420 433363 504476 433397
rect 504510 433363 504566 433397
rect 504600 433363 504774 433397
rect 504808 433363 504864 433397
rect 504898 433363 504954 433397
rect 504988 433363 505044 433397
rect 505078 433363 505134 433397
rect 505168 433363 505224 433397
rect 505258 433363 505314 433397
rect 505348 433363 505404 433397
rect 505438 433363 505494 433397
rect 505528 433363 505584 433397
rect 505618 433363 505674 433397
rect 505708 433363 505764 433397
rect 505798 433363 505854 433397
rect 505888 433363 506062 433397
rect 506096 433363 506152 433397
rect 506186 433363 506242 433397
rect 506276 433363 506332 433397
rect 506366 433363 506422 433397
rect 506456 433363 506512 433397
rect 506546 433363 506602 433397
rect 506636 433363 506692 433397
rect 506726 433363 506782 433397
rect 506816 433363 506872 433397
rect 506906 433363 506962 433397
rect 506996 433363 507052 433397
rect 507086 433363 507142 433397
rect 507176 433363 507350 433397
rect 507384 433363 507440 433397
rect 507474 433363 507530 433397
rect 507564 433363 507620 433397
rect 507654 433363 507710 433397
rect 507744 433363 507800 433397
rect 507834 433363 507890 433397
rect 507924 433363 507980 433397
rect 508014 433363 508070 433397
rect 508104 433363 508160 433397
rect 508194 433363 508250 433397
rect 508284 433363 508340 433397
rect 508374 433363 508430 433397
rect 508464 433363 508638 433397
rect 508672 433363 508728 433397
rect 508762 433363 508818 433397
rect 508852 433363 508908 433397
rect 508942 433363 508998 433397
rect 509032 433363 509088 433397
rect 509122 433363 509178 433397
rect 509212 433363 509268 433397
rect 509302 433363 509358 433397
rect 509392 433363 509448 433397
rect 509482 433363 509538 433397
rect 509572 433363 509628 433397
rect 509662 433363 509718 433397
rect 509752 433363 509926 433397
rect 509960 433363 510016 433397
rect 510050 433363 510106 433397
rect 510140 433363 510196 433397
rect 510230 433363 510286 433397
rect 510320 433363 510376 433397
rect 510410 433363 510466 433397
rect 510500 433363 510556 433397
rect 510590 433363 510646 433397
rect 510680 433363 510736 433397
rect 510770 433363 510826 433397
rect 510860 433363 510916 433397
rect 510950 433363 511006 433397
rect 511040 433363 511214 433397
rect 511248 433363 511304 433397
rect 511338 433363 511394 433397
rect 511428 433363 511484 433397
rect 511518 433363 511574 433397
rect 511608 433363 511664 433397
rect 511698 433363 511754 433397
rect 511788 433363 511844 433397
rect 511878 433363 511934 433397
rect 511968 433363 512024 433397
rect 512058 433363 512114 433397
rect 512148 433363 512204 433397
rect 512238 433363 512294 433397
rect 512328 433363 512502 433397
rect 512536 433363 512592 433397
rect 512626 433363 512682 433397
rect 512716 433363 512772 433397
rect 512806 433363 512862 433397
rect 512896 433363 512952 433397
rect 512986 433363 513042 433397
rect 513076 433363 513132 433397
rect 513166 433363 513222 433397
rect 513256 433363 513312 433397
rect 513346 433363 513402 433397
rect 513436 433363 513492 433397
rect 513526 433363 513582 433397
rect 513616 433363 513674 433397
rect 503370 433296 513674 433363
rect 503370 433262 503486 433296
rect 503520 433262 503576 433296
rect 503610 433262 503666 433296
rect 503700 433262 503756 433296
rect 503790 433262 503846 433296
rect 503880 433262 503936 433296
rect 503970 433262 504026 433296
rect 504060 433262 504116 433296
rect 504150 433262 504206 433296
rect 504240 433262 504296 433296
rect 504330 433262 504386 433296
rect 504420 433262 504476 433296
rect 504510 433262 504566 433296
rect 504600 433262 504774 433296
rect 504808 433262 504864 433296
rect 504898 433262 504954 433296
rect 504988 433262 505044 433296
rect 505078 433262 505134 433296
rect 505168 433262 505224 433296
rect 505258 433262 505314 433296
rect 505348 433262 505404 433296
rect 505438 433262 505494 433296
rect 505528 433262 505584 433296
rect 505618 433262 505674 433296
rect 505708 433262 505764 433296
rect 505798 433262 505854 433296
rect 505888 433262 506062 433296
rect 506096 433262 506152 433296
rect 506186 433262 506242 433296
rect 506276 433262 506332 433296
rect 506366 433262 506422 433296
rect 506456 433262 506512 433296
rect 506546 433262 506602 433296
rect 506636 433262 506692 433296
rect 506726 433262 506782 433296
rect 506816 433262 506872 433296
rect 506906 433262 506962 433296
rect 506996 433262 507052 433296
rect 507086 433262 507142 433296
rect 507176 433262 507350 433296
rect 507384 433262 507440 433296
rect 507474 433262 507530 433296
rect 507564 433262 507620 433296
rect 507654 433262 507710 433296
rect 507744 433262 507800 433296
rect 507834 433262 507890 433296
rect 507924 433262 507980 433296
rect 508014 433262 508070 433296
rect 508104 433262 508160 433296
rect 508194 433262 508250 433296
rect 508284 433262 508340 433296
rect 508374 433262 508430 433296
rect 508464 433262 508638 433296
rect 508672 433262 508728 433296
rect 508762 433262 508818 433296
rect 508852 433262 508908 433296
rect 508942 433262 508998 433296
rect 509032 433262 509088 433296
rect 509122 433262 509178 433296
rect 509212 433262 509268 433296
rect 509302 433262 509358 433296
rect 509392 433262 509448 433296
rect 509482 433262 509538 433296
rect 509572 433262 509628 433296
rect 509662 433262 509718 433296
rect 509752 433262 509926 433296
rect 509960 433262 510016 433296
rect 510050 433262 510106 433296
rect 510140 433262 510196 433296
rect 510230 433262 510286 433296
rect 510320 433262 510376 433296
rect 510410 433262 510466 433296
rect 510500 433262 510556 433296
rect 510590 433262 510646 433296
rect 510680 433262 510736 433296
rect 510770 433262 510826 433296
rect 510860 433262 510916 433296
rect 510950 433262 511006 433296
rect 511040 433262 511214 433296
rect 511248 433262 511304 433296
rect 511338 433262 511394 433296
rect 511428 433262 511484 433296
rect 511518 433262 511574 433296
rect 511608 433262 511664 433296
rect 511698 433262 511754 433296
rect 511788 433262 511844 433296
rect 511878 433262 511934 433296
rect 511968 433262 512024 433296
rect 512058 433262 512114 433296
rect 512148 433262 512204 433296
rect 512238 433262 512294 433296
rect 512328 433262 512502 433296
rect 512536 433262 512592 433296
rect 512626 433262 512682 433296
rect 512716 433262 512772 433296
rect 512806 433262 512862 433296
rect 512896 433262 512952 433296
rect 512986 433262 513042 433296
rect 513076 433262 513132 433296
rect 513166 433262 513222 433296
rect 513256 433262 513312 433296
rect 513346 433262 513402 433296
rect 513436 433262 513492 433296
rect 513526 433262 513582 433296
rect 513616 433262 513674 433296
rect 503370 433229 513674 433262
rect 503370 433200 503471 433229
rect 503370 433166 503402 433200
rect 503436 433166 503471 433200
rect 504557 433200 504759 433229
rect 503370 433110 503471 433166
rect 503370 433076 503402 433110
rect 503436 433076 503471 433110
rect 503370 433020 503471 433076
rect 503370 432986 503402 433020
rect 503436 432986 503471 433020
rect 503370 432930 503471 432986
rect 503370 432896 503402 432930
rect 503436 432896 503471 432930
rect 503370 432840 503471 432896
rect 503370 432806 503402 432840
rect 503436 432806 503471 432840
rect 503370 432750 503471 432806
rect 503370 432716 503402 432750
rect 503436 432716 503471 432750
rect 503370 432660 503471 432716
rect 503370 432626 503402 432660
rect 503436 432626 503471 432660
rect 503370 432570 503471 432626
rect 503370 432536 503402 432570
rect 503436 432536 503471 432570
rect 503370 432480 503471 432536
rect 503370 432446 503402 432480
rect 503436 432446 503471 432480
rect 503370 432390 503471 432446
rect 503370 432356 503402 432390
rect 503436 432356 503471 432390
rect 503370 432300 503471 432356
rect 503370 432266 503402 432300
rect 503436 432266 503471 432300
rect 503370 432210 503471 432266
rect 503370 432176 503402 432210
rect 503436 432176 503471 432210
rect 504557 433166 504589 433200
rect 504623 433166 504690 433200
rect 504724 433166 504759 433200
rect 505845 433200 506047 433229
rect 504557 433110 504759 433166
rect 504557 433076 504589 433110
rect 504623 433076 504690 433110
rect 504724 433076 504759 433110
rect 504557 433020 504759 433076
rect 504557 432986 504589 433020
rect 504623 432986 504690 433020
rect 504724 432986 504759 433020
rect 504557 432930 504759 432986
rect 504557 432896 504589 432930
rect 504623 432896 504690 432930
rect 504724 432896 504759 432930
rect 504557 432840 504759 432896
rect 504557 432806 504589 432840
rect 504623 432806 504690 432840
rect 504724 432806 504759 432840
rect 504557 432750 504759 432806
rect 504557 432716 504589 432750
rect 504623 432716 504690 432750
rect 504724 432716 504759 432750
rect 504557 432660 504759 432716
rect 504557 432626 504589 432660
rect 504623 432626 504690 432660
rect 504724 432626 504759 432660
rect 504557 432570 504759 432626
rect 504557 432536 504589 432570
rect 504623 432536 504690 432570
rect 504724 432536 504759 432570
rect 504557 432480 504759 432536
rect 504557 432446 504589 432480
rect 504623 432446 504690 432480
rect 504724 432446 504759 432480
rect 504557 432390 504759 432446
rect 504557 432356 504589 432390
rect 504623 432356 504690 432390
rect 504724 432356 504759 432390
rect 504557 432300 504759 432356
rect 504557 432266 504589 432300
rect 504623 432266 504690 432300
rect 504724 432266 504759 432300
rect 504557 432210 504759 432266
rect 503370 432143 503471 432176
rect 504557 432176 504589 432210
rect 504623 432176 504690 432210
rect 504724 432176 504759 432210
rect 505845 433166 505877 433200
rect 505911 433166 505978 433200
rect 506012 433166 506047 433200
rect 507133 433200 507335 433229
rect 505845 433110 506047 433166
rect 505845 433076 505877 433110
rect 505911 433076 505978 433110
rect 506012 433076 506047 433110
rect 505845 433020 506047 433076
rect 505845 432986 505877 433020
rect 505911 432986 505978 433020
rect 506012 432986 506047 433020
rect 505845 432930 506047 432986
rect 505845 432896 505877 432930
rect 505911 432896 505978 432930
rect 506012 432896 506047 432930
rect 505845 432840 506047 432896
rect 505845 432806 505877 432840
rect 505911 432806 505978 432840
rect 506012 432806 506047 432840
rect 505845 432750 506047 432806
rect 505845 432716 505877 432750
rect 505911 432716 505978 432750
rect 506012 432716 506047 432750
rect 505845 432660 506047 432716
rect 505845 432626 505877 432660
rect 505911 432626 505978 432660
rect 506012 432626 506047 432660
rect 505845 432570 506047 432626
rect 505845 432536 505877 432570
rect 505911 432536 505978 432570
rect 506012 432536 506047 432570
rect 505845 432480 506047 432536
rect 505845 432446 505877 432480
rect 505911 432446 505978 432480
rect 506012 432446 506047 432480
rect 505845 432390 506047 432446
rect 505845 432356 505877 432390
rect 505911 432356 505978 432390
rect 506012 432356 506047 432390
rect 505845 432300 506047 432356
rect 505845 432266 505877 432300
rect 505911 432266 505978 432300
rect 506012 432266 506047 432300
rect 505845 432210 506047 432266
rect 504557 432143 504759 432176
rect 505845 432176 505877 432210
rect 505911 432176 505978 432210
rect 506012 432176 506047 432210
rect 507133 433166 507165 433200
rect 507199 433166 507266 433200
rect 507300 433166 507335 433200
rect 508421 433200 508623 433229
rect 507133 433110 507335 433166
rect 507133 433076 507165 433110
rect 507199 433076 507266 433110
rect 507300 433076 507335 433110
rect 507133 433020 507335 433076
rect 507133 432986 507165 433020
rect 507199 432986 507266 433020
rect 507300 432986 507335 433020
rect 507133 432930 507335 432986
rect 507133 432896 507165 432930
rect 507199 432896 507266 432930
rect 507300 432896 507335 432930
rect 507133 432840 507335 432896
rect 507133 432806 507165 432840
rect 507199 432806 507266 432840
rect 507300 432806 507335 432840
rect 507133 432750 507335 432806
rect 507133 432716 507165 432750
rect 507199 432716 507266 432750
rect 507300 432716 507335 432750
rect 507133 432660 507335 432716
rect 507133 432626 507165 432660
rect 507199 432626 507266 432660
rect 507300 432626 507335 432660
rect 507133 432570 507335 432626
rect 507133 432536 507165 432570
rect 507199 432536 507266 432570
rect 507300 432536 507335 432570
rect 507133 432480 507335 432536
rect 507133 432446 507165 432480
rect 507199 432446 507266 432480
rect 507300 432446 507335 432480
rect 507133 432390 507335 432446
rect 507133 432356 507165 432390
rect 507199 432356 507266 432390
rect 507300 432356 507335 432390
rect 507133 432300 507335 432356
rect 507133 432266 507165 432300
rect 507199 432266 507266 432300
rect 507300 432266 507335 432300
rect 507133 432210 507335 432266
rect 505845 432143 506047 432176
rect 507133 432176 507165 432210
rect 507199 432176 507266 432210
rect 507300 432176 507335 432210
rect 508421 433166 508453 433200
rect 508487 433166 508554 433200
rect 508588 433166 508623 433200
rect 509709 433200 509911 433229
rect 508421 433110 508623 433166
rect 508421 433076 508453 433110
rect 508487 433076 508554 433110
rect 508588 433076 508623 433110
rect 508421 433020 508623 433076
rect 508421 432986 508453 433020
rect 508487 432986 508554 433020
rect 508588 432986 508623 433020
rect 508421 432930 508623 432986
rect 508421 432896 508453 432930
rect 508487 432896 508554 432930
rect 508588 432896 508623 432930
rect 508421 432840 508623 432896
rect 508421 432806 508453 432840
rect 508487 432806 508554 432840
rect 508588 432806 508623 432840
rect 508421 432750 508623 432806
rect 508421 432716 508453 432750
rect 508487 432716 508554 432750
rect 508588 432716 508623 432750
rect 508421 432660 508623 432716
rect 508421 432626 508453 432660
rect 508487 432626 508554 432660
rect 508588 432626 508623 432660
rect 508421 432570 508623 432626
rect 508421 432536 508453 432570
rect 508487 432536 508554 432570
rect 508588 432536 508623 432570
rect 508421 432480 508623 432536
rect 508421 432446 508453 432480
rect 508487 432446 508554 432480
rect 508588 432446 508623 432480
rect 508421 432390 508623 432446
rect 508421 432356 508453 432390
rect 508487 432356 508554 432390
rect 508588 432356 508623 432390
rect 508421 432300 508623 432356
rect 508421 432266 508453 432300
rect 508487 432266 508554 432300
rect 508588 432266 508623 432300
rect 508421 432210 508623 432266
rect 507133 432143 507335 432176
rect 508421 432176 508453 432210
rect 508487 432176 508554 432210
rect 508588 432176 508623 432210
rect 509709 433166 509741 433200
rect 509775 433166 509842 433200
rect 509876 433166 509911 433200
rect 510997 433200 511199 433229
rect 509709 433110 509911 433166
rect 509709 433076 509741 433110
rect 509775 433076 509842 433110
rect 509876 433076 509911 433110
rect 509709 433020 509911 433076
rect 509709 432986 509741 433020
rect 509775 432986 509842 433020
rect 509876 432986 509911 433020
rect 509709 432930 509911 432986
rect 509709 432896 509741 432930
rect 509775 432896 509842 432930
rect 509876 432896 509911 432930
rect 509709 432840 509911 432896
rect 509709 432806 509741 432840
rect 509775 432806 509842 432840
rect 509876 432806 509911 432840
rect 509709 432750 509911 432806
rect 509709 432716 509741 432750
rect 509775 432716 509842 432750
rect 509876 432716 509911 432750
rect 509709 432660 509911 432716
rect 509709 432626 509741 432660
rect 509775 432626 509842 432660
rect 509876 432626 509911 432660
rect 509709 432570 509911 432626
rect 509709 432536 509741 432570
rect 509775 432536 509842 432570
rect 509876 432536 509911 432570
rect 509709 432480 509911 432536
rect 509709 432446 509741 432480
rect 509775 432446 509842 432480
rect 509876 432446 509911 432480
rect 509709 432390 509911 432446
rect 509709 432356 509741 432390
rect 509775 432356 509842 432390
rect 509876 432356 509911 432390
rect 509709 432300 509911 432356
rect 509709 432266 509741 432300
rect 509775 432266 509842 432300
rect 509876 432266 509911 432300
rect 509709 432210 509911 432266
rect 508421 432143 508623 432176
rect 509709 432176 509741 432210
rect 509775 432176 509842 432210
rect 509876 432176 509911 432210
rect 510997 433166 511029 433200
rect 511063 433166 511130 433200
rect 511164 433166 511199 433200
rect 512285 433200 512487 433229
rect 510997 433110 511199 433166
rect 510997 433076 511029 433110
rect 511063 433076 511130 433110
rect 511164 433076 511199 433110
rect 510997 433020 511199 433076
rect 510997 432986 511029 433020
rect 511063 432986 511130 433020
rect 511164 432986 511199 433020
rect 510997 432930 511199 432986
rect 510997 432896 511029 432930
rect 511063 432896 511130 432930
rect 511164 432896 511199 432930
rect 510997 432840 511199 432896
rect 510997 432806 511029 432840
rect 511063 432806 511130 432840
rect 511164 432806 511199 432840
rect 510997 432750 511199 432806
rect 510997 432716 511029 432750
rect 511063 432716 511130 432750
rect 511164 432716 511199 432750
rect 510997 432660 511199 432716
rect 510997 432626 511029 432660
rect 511063 432626 511130 432660
rect 511164 432626 511199 432660
rect 510997 432570 511199 432626
rect 510997 432536 511029 432570
rect 511063 432536 511130 432570
rect 511164 432536 511199 432570
rect 510997 432480 511199 432536
rect 510997 432446 511029 432480
rect 511063 432446 511130 432480
rect 511164 432446 511199 432480
rect 510997 432390 511199 432446
rect 510997 432356 511029 432390
rect 511063 432356 511130 432390
rect 511164 432356 511199 432390
rect 510997 432300 511199 432356
rect 510997 432266 511029 432300
rect 511063 432266 511130 432300
rect 511164 432266 511199 432300
rect 510997 432210 511199 432266
rect 509709 432143 509911 432176
rect 510997 432176 511029 432210
rect 511063 432176 511130 432210
rect 511164 432176 511199 432210
rect 512285 433166 512317 433200
rect 512351 433166 512418 433200
rect 512452 433166 512487 433200
rect 513573 433200 513674 433229
rect 512285 433110 512487 433166
rect 512285 433076 512317 433110
rect 512351 433076 512418 433110
rect 512452 433076 512487 433110
rect 512285 433020 512487 433076
rect 512285 432986 512317 433020
rect 512351 432986 512418 433020
rect 512452 432986 512487 433020
rect 512285 432930 512487 432986
rect 512285 432896 512317 432930
rect 512351 432896 512418 432930
rect 512452 432896 512487 432930
rect 512285 432840 512487 432896
rect 512285 432806 512317 432840
rect 512351 432806 512418 432840
rect 512452 432806 512487 432840
rect 512285 432750 512487 432806
rect 512285 432716 512317 432750
rect 512351 432716 512418 432750
rect 512452 432716 512487 432750
rect 512285 432660 512487 432716
rect 512285 432626 512317 432660
rect 512351 432626 512418 432660
rect 512452 432626 512487 432660
rect 512285 432570 512487 432626
rect 512285 432536 512317 432570
rect 512351 432536 512418 432570
rect 512452 432536 512487 432570
rect 512285 432480 512487 432536
rect 512285 432446 512317 432480
rect 512351 432446 512418 432480
rect 512452 432446 512487 432480
rect 512285 432390 512487 432446
rect 512285 432356 512317 432390
rect 512351 432356 512418 432390
rect 512452 432356 512487 432390
rect 512285 432300 512487 432356
rect 512285 432266 512317 432300
rect 512351 432266 512418 432300
rect 512452 432266 512487 432300
rect 512285 432210 512487 432266
rect 510997 432143 511199 432176
rect 512285 432176 512317 432210
rect 512351 432176 512418 432210
rect 512452 432176 512487 432210
rect 513573 433166 513605 433200
rect 513639 433166 513674 433200
rect 513573 433110 513674 433166
rect 513573 433076 513605 433110
rect 513639 433076 513674 433110
rect 513573 433020 513674 433076
rect 513573 432986 513605 433020
rect 513639 432986 513674 433020
rect 513573 432930 513674 432986
rect 513573 432896 513605 432930
rect 513639 432896 513674 432930
rect 513573 432840 513674 432896
rect 513573 432806 513605 432840
rect 513639 432806 513674 432840
rect 513573 432750 513674 432806
rect 513573 432716 513605 432750
rect 513639 432716 513674 432750
rect 513573 432660 513674 432716
rect 513573 432626 513605 432660
rect 513639 432626 513674 432660
rect 513573 432570 513674 432626
rect 513573 432536 513605 432570
rect 513639 432536 513674 432570
rect 513573 432480 513674 432536
rect 513573 432446 513605 432480
rect 513639 432446 513674 432480
rect 513573 432390 513674 432446
rect 513573 432356 513605 432390
rect 513639 432356 513674 432390
rect 513573 432300 513674 432356
rect 513573 432266 513605 432300
rect 513639 432266 513674 432300
rect 513573 432210 513674 432266
rect 512285 432143 512487 432176
rect 513573 432176 513605 432210
rect 513639 432176 513674 432210
rect 513573 432143 513674 432176
rect 503370 432109 513674 432143
rect 503370 432075 503486 432109
rect 503520 432075 503576 432109
rect 503610 432075 503666 432109
rect 503700 432075 503756 432109
rect 503790 432075 503846 432109
rect 503880 432075 503936 432109
rect 503970 432075 504026 432109
rect 504060 432075 504116 432109
rect 504150 432075 504206 432109
rect 504240 432075 504296 432109
rect 504330 432075 504386 432109
rect 504420 432075 504476 432109
rect 504510 432075 504566 432109
rect 504600 432075 504774 432109
rect 504808 432075 504864 432109
rect 504898 432075 504954 432109
rect 504988 432075 505044 432109
rect 505078 432075 505134 432109
rect 505168 432075 505224 432109
rect 505258 432075 505314 432109
rect 505348 432075 505404 432109
rect 505438 432075 505494 432109
rect 505528 432075 505584 432109
rect 505618 432075 505674 432109
rect 505708 432075 505764 432109
rect 505798 432075 505854 432109
rect 505888 432075 506062 432109
rect 506096 432075 506152 432109
rect 506186 432075 506242 432109
rect 506276 432075 506332 432109
rect 506366 432075 506422 432109
rect 506456 432075 506512 432109
rect 506546 432075 506602 432109
rect 506636 432075 506692 432109
rect 506726 432075 506782 432109
rect 506816 432075 506872 432109
rect 506906 432075 506962 432109
rect 506996 432075 507052 432109
rect 507086 432075 507142 432109
rect 507176 432075 507350 432109
rect 507384 432075 507440 432109
rect 507474 432075 507530 432109
rect 507564 432075 507620 432109
rect 507654 432075 507710 432109
rect 507744 432075 507800 432109
rect 507834 432075 507890 432109
rect 507924 432075 507980 432109
rect 508014 432075 508070 432109
rect 508104 432075 508160 432109
rect 508194 432075 508250 432109
rect 508284 432075 508340 432109
rect 508374 432075 508430 432109
rect 508464 432075 508638 432109
rect 508672 432075 508728 432109
rect 508762 432075 508818 432109
rect 508852 432075 508908 432109
rect 508942 432075 508998 432109
rect 509032 432075 509088 432109
rect 509122 432075 509178 432109
rect 509212 432075 509268 432109
rect 509302 432075 509358 432109
rect 509392 432075 509448 432109
rect 509482 432075 509538 432109
rect 509572 432075 509628 432109
rect 509662 432075 509718 432109
rect 509752 432075 509926 432109
rect 509960 432075 510016 432109
rect 510050 432075 510106 432109
rect 510140 432075 510196 432109
rect 510230 432075 510286 432109
rect 510320 432075 510376 432109
rect 510410 432075 510466 432109
rect 510500 432075 510556 432109
rect 510590 432075 510646 432109
rect 510680 432075 510736 432109
rect 510770 432075 510826 432109
rect 510860 432075 510916 432109
rect 510950 432075 511006 432109
rect 511040 432075 511214 432109
rect 511248 432075 511304 432109
rect 511338 432075 511394 432109
rect 511428 432075 511484 432109
rect 511518 432075 511574 432109
rect 511608 432075 511664 432109
rect 511698 432075 511754 432109
rect 511788 432075 511844 432109
rect 511878 432075 511934 432109
rect 511968 432075 512024 432109
rect 512058 432075 512114 432109
rect 512148 432075 512204 432109
rect 512238 432075 512294 432109
rect 512328 432075 512502 432109
rect 512536 432075 512592 432109
rect 512626 432075 512682 432109
rect 512716 432075 512772 432109
rect 512806 432075 512862 432109
rect 512896 432075 512952 432109
rect 512986 432075 513042 432109
rect 513076 432075 513132 432109
rect 513166 432075 513222 432109
rect 513256 432075 513312 432109
rect 513346 432075 513402 432109
rect 513436 432075 513492 432109
rect 513526 432075 513582 432109
rect 513616 432075 513674 432109
rect 503370 431068 513674 432075
rect 500320 431044 526592 431068
rect 500320 430044 500344 431044
rect 526568 430044 526592 431044
rect 500320 430020 526592 430044
rect 527568 430020 527592 475332
rect 528592 430020 528616 475332
rect 572316 455212 572412 455246
rect 577642 455212 577738 455246
rect 572316 455150 572350 455212
rect 577704 455150 577738 455212
rect 572316 453994 572350 454056
rect 577704 453994 577738 454056
rect 572316 453960 572412 453994
rect 577642 453960 577738 453994
rect 527568 429996 528616 430020
<< nsubdiff >>
rect 562156 495480 562252 495514
rect 567482 495480 567578 495514
rect 562156 495417 562190 495480
rect 567544 495417 567578 495480
rect 562156 494252 562190 494315
rect 567544 494252 567578 494315
rect 562156 494218 562252 494252
rect 567482 494218 567578 494252
rect 503126 470202 505668 470252
rect 503126 470102 503226 470202
rect 505568 470102 505668 470202
rect 503126 470052 505668 470102
rect 502572 466620 502772 466720
rect 502572 464278 502622 466620
rect 502722 464278 502772 466620
rect 502572 464178 502772 464278
rect 503126 461074 505668 461124
rect 503126 460974 503226 461074
rect 505568 460974 505668 461074
rect 503126 460924 505668 460974
rect 503328 460252 510728 460452
rect 503328 460052 503528 460252
rect 510528 460052 510728 460252
rect 503328 459852 510728 460052
rect 503328 454342 510728 454542
rect 503328 454142 503528 454342
rect 510528 454142 510728 454342
rect 503328 453942 510728 454142
rect 503328 448842 510728 449042
rect 503328 448642 503528 448842
rect 510528 448642 510728 448842
rect 503328 448442 510728 448642
rect 503326 442886 510726 443086
rect 503326 442686 503526 442886
rect 510526 442686 510726 442886
rect 503326 442486 510726 442686
rect 503533 438300 504495 438319
rect 503533 438266 503665 438300
rect 503699 438266 503755 438300
rect 503789 438266 503845 438300
rect 503879 438266 503935 438300
rect 503969 438266 504025 438300
rect 504059 438266 504115 438300
rect 504149 438266 504205 438300
rect 504239 438266 504295 438300
rect 504329 438266 504385 438300
rect 504419 438266 504495 438300
rect 503533 438247 504495 438266
rect 503533 438222 503605 438247
rect 503533 438188 503552 438222
rect 503586 438188 503605 438222
rect 503533 438132 503605 438188
rect 504423 438188 504495 438247
rect 503533 438098 503552 438132
rect 503586 438098 503605 438132
rect 503533 438042 503605 438098
rect 503533 438008 503552 438042
rect 503586 438008 503605 438042
rect 503533 437952 503605 438008
rect 503533 437918 503552 437952
rect 503586 437918 503605 437952
rect 503533 437862 503605 437918
rect 503533 437828 503552 437862
rect 503586 437828 503605 437862
rect 503533 437772 503605 437828
rect 503533 437738 503552 437772
rect 503586 437738 503605 437772
rect 503533 437682 503605 437738
rect 503533 437648 503552 437682
rect 503586 437648 503605 437682
rect 503533 437592 503605 437648
rect 503533 437558 503552 437592
rect 503586 437558 503605 437592
rect 503533 437502 503605 437558
rect 503533 437468 503552 437502
rect 503586 437468 503605 437502
rect 504423 438154 504442 438188
rect 504476 438154 504495 438188
rect 504423 438098 504495 438154
rect 504423 438064 504442 438098
rect 504476 438064 504495 438098
rect 504423 438008 504495 438064
rect 504423 437974 504442 438008
rect 504476 437974 504495 438008
rect 504423 437918 504495 437974
rect 504423 437884 504442 437918
rect 504476 437884 504495 437918
rect 504423 437828 504495 437884
rect 504423 437794 504442 437828
rect 504476 437794 504495 437828
rect 504423 437738 504495 437794
rect 504423 437704 504442 437738
rect 504476 437704 504495 437738
rect 504423 437648 504495 437704
rect 504423 437614 504442 437648
rect 504476 437614 504495 437648
rect 504423 437558 504495 437614
rect 504423 437524 504442 437558
rect 504476 437524 504495 437558
rect 503533 437429 503605 437468
rect 504423 437468 504495 437524
rect 504423 437434 504442 437468
rect 504476 437434 504495 437468
rect 504423 437429 504495 437434
rect 503533 437410 504495 437429
rect 503533 437376 503646 437410
rect 503680 437376 503736 437410
rect 503770 437376 503826 437410
rect 503860 437376 503916 437410
rect 503950 437376 504006 437410
rect 504040 437376 504096 437410
rect 504130 437376 504186 437410
rect 504220 437376 504276 437410
rect 504310 437376 504366 437410
rect 504400 437376 504495 437410
rect 503533 437357 504495 437376
rect 504821 438300 505783 438319
rect 504821 438266 504953 438300
rect 504987 438266 505043 438300
rect 505077 438266 505133 438300
rect 505167 438266 505223 438300
rect 505257 438266 505313 438300
rect 505347 438266 505403 438300
rect 505437 438266 505493 438300
rect 505527 438266 505583 438300
rect 505617 438266 505673 438300
rect 505707 438266 505783 438300
rect 504821 438247 505783 438266
rect 504821 438222 504893 438247
rect 504821 438188 504840 438222
rect 504874 438188 504893 438222
rect 504821 438132 504893 438188
rect 505711 438188 505783 438247
rect 504821 438098 504840 438132
rect 504874 438098 504893 438132
rect 504821 438042 504893 438098
rect 504821 438008 504840 438042
rect 504874 438008 504893 438042
rect 504821 437952 504893 438008
rect 504821 437918 504840 437952
rect 504874 437918 504893 437952
rect 504821 437862 504893 437918
rect 504821 437828 504840 437862
rect 504874 437828 504893 437862
rect 504821 437772 504893 437828
rect 504821 437738 504840 437772
rect 504874 437738 504893 437772
rect 504821 437682 504893 437738
rect 504821 437648 504840 437682
rect 504874 437648 504893 437682
rect 504821 437592 504893 437648
rect 504821 437558 504840 437592
rect 504874 437558 504893 437592
rect 504821 437502 504893 437558
rect 504821 437468 504840 437502
rect 504874 437468 504893 437502
rect 505711 438154 505730 438188
rect 505764 438154 505783 438188
rect 505711 438098 505783 438154
rect 505711 438064 505730 438098
rect 505764 438064 505783 438098
rect 505711 438008 505783 438064
rect 505711 437974 505730 438008
rect 505764 437974 505783 438008
rect 505711 437918 505783 437974
rect 505711 437884 505730 437918
rect 505764 437884 505783 437918
rect 505711 437828 505783 437884
rect 505711 437794 505730 437828
rect 505764 437794 505783 437828
rect 505711 437738 505783 437794
rect 505711 437704 505730 437738
rect 505764 437704 505783 437738
rect 505711 437648 505783 437704
rect 505711 437614 505730 437648
rect 505764 437614 505783 437648
rect 505711 437558 505783 437614
rect 505711 437524 505730 437558
rect 505764 437524 505783 437558
rect 504821 437429 504893 437468
rect 505711 437468 505783 437524
rect 505711 437434 505730 437468
rect 505764 437434 505783 437468
rect 505711 437429 505783 437434
rect 504821 437410 505783 437429
rect 504821 437376 504934 437410
rect 504968 437376 505024 437410
rect 505058 437376 505114 437410
rect 505148 437376 505204 437410
rect 505238 437376 505294 437410
rect 505328 437376 505384 437410
rect 505418 437376 505474 437410
rect 505508 437376 505564 437410
rect 505598 437376 505654 437410
rect 505688 437376 505783 437410
rect 504821 437357 505783 437376
rect 506109 438300 507071 438319
rect 506109 438266 506241 438300
rect 506275 438266 506331 438300
rect 506365 438266 506421 438300
rect 506455 438266 506511 438300
rect 506545 438266 506601 438300
rect 506635 438266 506691 438300
rect 506725 438266 506781 438300
rect 506815 438266 506871 438300
rect 506905 438266 506961 438300
rect 506995 438266 507071 438300
rect 506109 438247 507071 438266
rect 506109 438222 506181 438247
rect 506109 438188 506128 438222
rect 506162 438188 506181 438222
rect 506109 438132 506181 438188
rect 506999 438188 507071 438247
rect 506109 438098 506128 438132
rect 506162 438098 506181 438132
rect 506109 438042 506181 438098
rect 506109 438008 506128 438042
rect 506162 438008 506181 438042
rect 506109 437952 506181 438008
rect 506109 437918 506128 437952
rect 506162 437918 506181 437952
rect 506109 437862 506181 437918
rect 506109 437828 506128 437862
rect 506162 437828 506181 437862
rect 506109 437772 506181 437828
rect 506109 437738 506128 437772
rect 506162 437738 506181 437772
rect 506109 437682 506181 437738
rect 506109 437648 506128 437682
rect 506162 437648 506181 437682
rect 506109 437592 506181 437648
rect 506109 437558 506128 437592
rect 506162 437558 506181 437592
rect 506109 437502 506181 437558
rect 506109 437468 506128 437502
rect 506162 437468 506181 437502
rect 506999 438154 507018 438188
rect 507052 438154 507071 438188
rect 506999 438098 507071 438154
rect 506999 438064 507018 438098
rect 507052 438064 507071 438098
rect 506999 438008 507071 438064
rect 506999 437974 507018 438008
rect 507052 437974 507071 438008
rect 506999 437918 507071 437974
rect 506999 437884 507018 437918
rect 507052 437884 507071 437918
rect 506999 437828 507071 437884
rect 506999 437794 507018 437828
rect 507052 437794 507071 437828
rect 506999 437738 507071 437794
rect 506999 437704 507018 437738
rect 507052 437704 507071 437738
rect 506999 437648 507071 437704
rect 506999 437614 507018 437648
rect 507052 437614 507071 437648
rect 506999 437558 507071 437614
rect 506999 437524 507018 437558
rect 507052 437524 507071 437558
rect 506109 437429 506181 437468
rect 506999 437468 507071 437524
rect 506999 437434 507018 437468
rect 507052 437434 507071 437468
rect 506999 437429 507071 437434
rect 506109 437410 507071 437429
rect 506109 437376 506222 437410
rect 506256 437376 506312 437410
rect 506346 437376 506402 437410
rect 506436 437376 506492 437410
rect 506526 437376 506582 437410
rect 506616 437376 506672 437410
rect 506706 437376 506762 437410
rect 506796 437376 506852 437410
rect 506886 437376 506942 437410
rect 506976 437376 507071 437410
rect 506109 437357 507071 437376
rect 507397 438300 508359 438319
rect 507397 438266 507529 438300
rect 507563 438266 507619 438300
rect 507653 438266 507709 438300
rect 507743 438266 507799 438300
rect 507833 438266 507889 438300
rect 507923 438266 507979 438300
rect 508013 438266 508069 438300
rect 508103 438266 508159 438300
rect 508193 438266 508249 438300
rect 508283 438266 508359 438300
rect 507397 438247 508359 438266
rect 507397 438222 507469 438247
rect 507397 438188 507416 438222
rect 507450 438188 507469 438222
rect 507397 438132 507469 438188
rect 508287 438188 508359 438247
rect 507397 438098 507416 438132
rect 507450 438098 507469 438132
rect 507397 438042 507469 438098
rect 507397 438008 507416 438042
rect 507450 438008 507469 438042
rect 507397 437952 507469 438008
rect 507397 437918 507416 437952
rect 507450 437918 507469 437952
rect 507397 437862 507469 437918
rect 507397 437828 507416 437862
rect 507450 437828 507469 437862
rect 507397 437772 507469 437828
rect 507397 437738 507416 437772
rect 507450 437738 507469 437772
rect 507397 437682 507469 437738
rect 507397 437648 507416 437682
rect 507450 437648 507469 437682
rect 507397 437592 507469 437648
rect 507397 437558 507416 437592
rect 507450 437558 507469 437592
rect 507397 437502 507469 437558
rect 507397 437468 507416 437502
rect 507450 437468 507469 437502
rect 508287 438154 508306 438188
rect 508340 438154 508359 438188
rect 508287 438098 508359 438154
rect 508287 438064 508306 438098
rect 508340 438064 508359 438098
rect 508287 438008 508359 438064
rect 508287 437974 508306 438008
rect 508340 437974 508359 438008
rect 508287 437918 508359 437974
rect 508287 437884 508306 437918
rect 508340 437884 508359 437918
rect 508287 437828 508359 437884
rect 508287 437794 508306 437828
rect 508340 437794 508359 437828
rect 508287 437738 508359 437794
rect 508287 437704 508306 437738
rect 508340 437704 508359 437738
rect 508287 437648 508359 437704
rect 508287 437614 508306 437648
rect 508340 437614 508359 437648
rect 508287 437558 508359 437614
rect 508287 437524 508306 437558
rect 508340 437524 508359 437558
rect 507397 437429 507469 437468
rect 508287 437468 508359 437524
rect 508287 437434 508306 437468
rect 508340 437434 508359 437468
rect 508287 437429 508359 437434
rect 507397 437410 508359 437429
rect 507397 437376 507510 437410
rect 507544 437376 507600 437410
rect 507634 437376 507690 437410
rect 507724 437376 507780 437410
rect 507814 437376 507870 437410
rect 507904 437376 507960 437410
rect 507994 437376 508050 437410
rect 508084 437376 508140 437410
rect 508174 437376 508230 437410
rect 508264 437376 508359 437410
rect 507397 437357 508359 437376
rect 508685 438300 509647 438319
rect 508685 438266 508817 438300
rect 508851 438266 508907 438300
rect 508941 438266 508997 438300
rect 509031 438266 509087 438300
rect 509121 438266 509177 438300
rect 509211 438266 509267 438300
rect 509301 438266 509357 438300
rect 509391 438266 509447 438300
rect 509481 438266 509537 438300
rect 509571 438266 509647 438300
rect 508685 438247 509647 438266
rect 508685 438222 508757 438247
rect 508685 438188 508704 438222
rect 508738 438188 508757 438222
rect 508685 438132 508757 438188
rect 509575 438188 509647 438247
rect 508685 438098 508704 438132
rect 508738 438098 508757 438132
rect 508685 438042 508757 438098
rect 508685 438008 508704 438042
rect 508738 438008 508757 438042
rect 508685 437952 508757 438008
rect 508685 437918 508704 437952
rect 508738 437918 508757 437952
rect 508685 437862 508757 437918
rect 508685 437828 508704 437862
rect 508738 437828 508757 437862
rect 508685 437772 508757 437828
rect 508685 437738 508704 437772
rect 508738 437738 508757 437772
rect 508685 437682 508757 437738
rect 508685 437648 508704 437682
rect 508738 437648 508757 437682
rect 508685 437592 508757 437648
rect 508685 437558 508704 437592
rect 508738 437558 508757 437592
rect 508685 437502 508757 437558
rect 508685 437468 508704 437502
rect 508738 437468 508757 437502
rect 509575 438154 509594 438188
rect 509628 438154 509647 438188
rect 509575 438098 509647 438154
rect 509575 438064 509594 438098
rect 509628 438064 509647 438098
rect 509575 438008 509647 438064
rect 509575 437974 509594 438008
rect 509628 437974 509647 438008
rect 509575 437918 509647 437974
rect 509575 437884 509594 437918
rect 509628 437884 509647 437918
rect 509575 437828 509647 437884
rect 509575 437794 509594 437828
rect 509628 437794 509647 437828
rect 509575 437738 509647 437794
rect 509575 437704 509594 437738
rect 509628 437704 509647 437738
rect 509575 437648 509647 437704
rect 509575 437614 509594 437648
rect 509628 437614 509647 437648
rect 509575 437558 509647 437614
rect 509575 437524 509594 437558
rect 509628 437524 509647 437558
rect 508685 437429 508757 437468
rect 509575 437468 509647 437524
rect 509575 437434 509594 437468
rect 509628 437434 509647 437468
rect 509575 437429 509647 437434
rect 508685 437410 509647 437429
rect 508685 437376 508798 437410
rect 508832 437376 508888 437410
rect 508922 437376 508978 437410
rect 509012 437376 509068 437410
rect 509102 437376 509158 437410
rect 509192 437376 509248 437410
rect 509282 437376 509338 437410
rect 509372 437376 509428 437410
rect 509462 437376 509518 437410
rect 509552 437376 509647 437410
rect 508685 437357 509647 437376
rect 509973 438300 510935 438319
rect 509973 438266 510105 438300
rect 510139 438266 510195 438300
rect 510229 438266 510285 438300
rect 510319 438266 510375 438300
rect 510409 438266 510465 438300
rect 510499 438266 510555 438300
rect 510589 438266 510645 438300
rect 510679 438266 510735 438300
rect 510769 438266 510825 438300
rect 510859 438266 510935 438300
rect 509973 438247 510935 438266
rect 509973 438222 510045 438247
rect 509973 438188 509992 438222
rect 510026 438188 510045 438222
rect 509973 438132 510045 438188
rect 510863 438188 510935 438247
rect 509973 438098 509992 438132
rect 510026 438098 510045 438132
rect 509973 438042 510045 438098
rect 509973 438008 509992 438042
rect 510026 438008 510045 438042
rect 509973 437952 510045 438008
rect 509973 437918 509992 437952
rect 510026 437918 510045 437952
rect 509973 437862 510045 437918
rect 509973 437828 509992 437862
rect 510026 437828 510045 437862
rect 509973 437772 510045 437828
rect 509973 437738 509992 437772
rect 510026 437738 510045 437772
rect 509973 437682 510045 437738
rect 509973 437648 509992 437682
rect 510026 437648 510045 437682
rect 509973 437592 510045 437648
rect 509973 437558 509992 437592
rect 510026 437558 510045 437592
rect 509973 437502 510045 437558
rect 509973 437468 509992 437502
rect 510026 437468 510045 437502
rect 510863 438154 510882 438188
rect 510916 438154 510935 438188
rect 510863 438098 510935 438154
rect 510863 438064 510882 438098
rect 510916 438064 510935 438098
rect 510863 438008 510935 438064
rect 510863 437974 510882 438008
rect 510916 437974 510935 438008
rect 510863 437918 510935 437974
rect 510863 437884 510882 437918
rect 510916 437884 510935 437918
rect 510863 437828 510935 437884
rect 510863 437794 510882 437828
rect 510916 437794 510935 437828
rect 510863 437738 510935 437794
rect 510863 437704 510882 437738
rect 510916 437704 510935 437738
rect 510863 437648 510935 437704
rect 510863 437614 510882 437648
rect 510916 437614 510935 437648
rect 510863 437558 510935 437614
rect 510863 437524 510882 437558
rect 510916 437524 510935 437558
rect 509973 437429 510045 437468
rect 510863 437468 510935 437524
rect 510863 437434 510882 437468
rect 510916 437434 510935 437468
rect 510863 437429 510935 437434
rect 509973 437410 510935 437429
rect 509973 437376 510086 437410
rect 510120 437376 510176 437410
rect 510210 437376 510266 437410
rect 510300 437376 510356 437410
rect 510390 437376 510446 437410
rect 510480 437376 510536 437410
rect 510570 437376 510626 437410
rect 510660 437376 510716 437410
rect 510750 437376 510806 437410
rect 510840 437376 510935 437410
rect 509973 437357 510935 437376
rect 511261 438300 512223 438319
rect 511261 438266 511393 438300
rect 511427 438266 511483 438300
rect 511517 438266 511573 438300
rect 511607 438266 511663 438300
rect 511697 438266 511753 438300
rect 511787 438266 511843 438300
rect 511877 438266 511933 438300
rect 511967 438266 512023 438300
rect 512057 438266 512113 438300
rect 512147 438266 512223 438300
rect 511261 438247 512223 438266
rect 511261 438222 511333 438247
rect 511261 438188 511280 438222
rect 511314 438188 511333 438222
rect 511261 438132 511333 438188
rect 512151 438188 512223 438247
rect 511261 438098 511280 438132
rect 511314 438098 511333 438132
rect 511261 438042 511333 438098
rect 511261 438008 511280 438042
rect 511314 438008 511333 438042
rect 511261 437952 511333 438008
rect 511261 437918 511280 437952
rect 511314 437918 511333 437952
rect 511261 437862 511333 437918
rect 511261 437828 511280 437862
rect 511314 437828 511333 437862
rect 511261 437772 511333 437828
rect 511261 437738 511280 437772
rect 511314 437738 511333 437772
rect 511261 437682 511333 437738
rect 511261 437648 511280 437682
rect 511314 437648 511333 437682
rect 511261 437592 511333 437648
rect 511261 437558 511280 437592
rect 511314 437558 511333 437592
rect 511261 437502 511333 437558
rect 511261 437468 511280 437502
rect 511314 437468 511333 437502
rect 512151 438154 512170 438188
rect 512204 438154 512223 438188
rect 512151 438098 512223 438154
rect 512151 438064 512170 438098
rect 512204 438064 512223 438098
rect 512151 438008 512223 438064
rect 512151 437974 512170 438008
rect 512204 437974 512223 438008
rect 512151 437918 512223 437974
rect 512151 437884 512170 437918
rect 512204 437884 512223 437918
rect 512151 437828 512223 437884
rect 512151 437794 512170 437828
rect 512204 437794 512223 437828
rect 512151 437738 512223 437794
rect 512151 437704 512170 437738
rect 512204 437704 512223 437738
rect 512151 437648 512223 437704
rect 512151 437614 512170 437648
rect 512204 437614 512223 437648
rect 512151 437558 512223 437614
rect 512151 437524 512170 437558
rect 512204 437524 512223 437558
rect 511261 437429 511333 437468
rect 512151 437468 512223 437524
rect 512151 437434 512170 437468
rect 512204 437434 512223 437468
rect 512151 437429 512223 437434
rect 511261 437410 512223 437429
rect 511261 437376 511374 437410
rect 511408 437376 511464 437410
rect 511498 437376 511554 437410
rect 511588 437376 511644 437410
rect 511678 437376 511734 437410
rect 511768 437376 511824 437410
rect 511858 437376 511914 437410
rect 511948 437376 512004 437410
rect 512038 437376 512094 437410
rect 512128 437376 512223 437410
rect 511261 437357 512223 437376
rect 512549 438300 513511 438319
rect 512549 438266 512681 438300
rect 512715 438266 512771 438300
rect 512805 438266 512861 438300
rect 512895 438266 512951 438300
rect 512985 438266 513041 438300
rect 513075 438266 513131 438300
rect 513165 438266 513221 438300
rect 513255 438266 513311 438300
rect 513345 438266 513401 438300
rect 513435 438266 513511 438300
rect 512549 438247 513511 438266
rect 512549 438222 512621 438247
rect 512549 438188 512568 438222
rect 512602 438188 512621 438222
rect 512549 438132 512621 438188
rect 513439 438188 513511 438247
rect 512549 438098 512568 438132
rect 512602 438098 512621 438132
rect 512549 438042 512621 438098
rect 512549 438008 512568 438042
rect 512602 438008 512621 438042
rect 512549 437952 512621 438008
rect 512549 437918 512568 437952
rect 512602 437918 512621 437952
rect 512549 437862 512621 437918
rect 512549 437828 512568 437862
rect 512602 437828 512621 437862
rect 512549 437772 512621 437828
rect 512549 437738 512568 437772
rect 512602 437738 512621 437772
rect 512549 437682 512621 437738
rect 512549 437648 512568 437682
rect 512602 437648 512621 437682
rect 512549 437592 512621 437648
rect 512549 437558 512568 437592
rect 512602 437558 512621 437592
rect 512549 437502 512621 437558
rect 512549 437468 512568 437502
rect 512602 437468 512621 437502
rect 513439 438154 513458 438188
rect 513492 438154 513511 438188
rect 513439 438098 513511 438154
rect 513439 438064 513458 438098
rect 513492 438064 513511 438098
rect 513439 438008 513511 438064
rect 513439 437974 513458 438008
rect 513492 437974 513511 438008
rect 513439 437918 513511 437974
rect 513439 437884 513458 437918
rect 513492 437884 513511 437918
rect 513439 437828 513511 437884
rect 513439 437794 513458 437828
rect 513492 437794 513511 437828
rect 513439 437738 513511 437794
rect 513439 437704 513458 437738
rect 513492 437704 513511 437738
rect 513439 437648 513511 437704
rect 513439 437614 513458 437648
rect 513492 437614 513511 437648
rect 513439 437558 513511 437614
rect 513439 437524 513458 437558
rect 513492 437524 513511 437558
rect 512549 437429 512621 437468
rect 513439 437468 513511 437524
rect 513439 437434 513458 437468
rect 513492 437434 513511 437468
rect 513439 437429 513511 437434
rect 512549 437410 513511 437429
rect 512549 437376 512662 437410
rect 512696 437376 512752 437410
rect 512786 437376 512842 437410
rect 512876 437376 512932 437410
rect 512966 437376 513022 437410
rect 513056 437376 513112 437410
rect 513146 437376 513202 437410
rect 513236 437376 513292 437410
rect 513326 437376 513382 437410
rect 513416 437376 513511 437410
rect 512549 437357 513511 437376
rect 503533 437012 504495 437031
rect 503533 436978 503665 437012
rect 503699 436978 503755 437012
rect 503789 436978 503845 437012
rect 503879 436978 503935 437012
rect 503969 436978 504025 437012
rect 504059 436978 504115 437012
rect 504149 436978 504205 437012
rect 504239 436978 504295 437012
rect 504329 436978 504385 437012
rect 504419 436978 504495 437012
rect 503533 436959 504495 436978
rect 503533 436934 503605 436959
rect 503533 436900 503552 436934
rect 503586 436900 503605 436934
rect 503533 436844 503605 436900
rect 504423 436900 504495 436959
rect 503533 436810 503552 436844
rect 503586 436810 503605 436844
rect 503533 436754 503605 436810
rect 503533 436720 503552 436754
rect 503586 436720 503605 436754
rect 503533 436664 503605 436720
rect 503533 436630 503552 436664
rect 503586 436630 503605 436664
rect 503533 436574 503605 436630
rect 503533 436540 503552 436574
rect 503586 436540 503605 436574
rect 503533 436484 503605 436540
rect 503533 436450 503552 436484
rect 503586 436450 503605 436484
rect 503533 436394 503605 436450
rect 503533 436360 503552 436394
rect 503586 436360 503605 436394
rect 503533 436304 503605 436360
rect 503533 436270 503552 436304
rect 503586 436270 503605 436304
rect 503533 436214 503605 436270
rect 503533 436180 503552 436214
rect 503586 436180 503605 436214
rect 504423 436866 504442 436900
rect 504476 436866 504495 436900
rect 504423 436810 504495 436866
rect 504423 436776 504442 436810
rect 504476 436776 504495 436810
rect 504423 436720 504495 436776
rect 504423 436686 504442 436720
rect 504476 436686 504495 436720
rect 504423 436630 504495 436686
rect 504423 436596 504442 436630
rect 504476 436596 504495 436630
rect 504423 436540 504495 436596
rect 504423 436506 504442 436540
rect 504476 436506 504495 436540
rect 504423 436450 504495 436506
rect 504423 436416 504442 436450
rect 504476 436416 504495 436450
rect 504423 436360 504495 436416
rect 504423 436326 504442 436360
rect 504476 436326 504495 436360
rect 504423 436270 504495 436326
rect 504423 436236 504442 436270
rect 504476 436236 504495 436270
rect 503533 436141 503605 436180
rect 504423 436180 504495 436236
rect 504423 436146 504442 436180
rect 504476 436146 504495 436180
rect 504423 436141 504495 436146
rect 503533 436122 504495 436141
rect 503533 436088 503646 436122
rect 503680 436088 503736 436122
rect 503770 436088 503826 436122
rect 503860 436088 503916 436122
rect 503950 436088 504006 436122
rect 504040 436088 504096 436122
rect 504130 436088 504186 436122
rect 504220 436088 504276 436122
rect 504310 436088 504366 436122
rect 504400 436088 504495 436122
rect 503533 436069 504495 436088
rect 504821 437012 505783 437031
rect 504821 436978 504953 437012
rect 504987 436978 505043 437012
rect 505077 436978 505133 437012
rect 505167 436978 505223 437012
rect 505257 436978 505313 437012
rect 505347 436978 505403 437012
rect 505437 436978 505493 437012
rect 505527 436978 505583 437012
rect 505617 436978 505673 437012
rect 505707 436978 505783 437012
rect 504821 436959 505783 436978
rect 504821 436934 504893 436959
rect 504821 436900 504840 436934
rect 504874 436900 504893 436934
rect 504821 436844 504893 436900
rect 505711 436900 505783 436959
rect 504821 436810 504840 436844
rect 504874 436810 504893 436844
rect 504821 436754 504893 436810
rect 504821 436720 504840 436754
rect 504874 436720 504893 436754
rect 504821 436664 504893 436720
rect 504821 436630 504840 436664
rect 504874 436630 504893 436664
rect 504821 436574 504893 436630
rect 504821 436540 504840 436574
rect 504874 436540 504893 436574
rect 504821 436484 504893 436540
rect 504821 436450 504840 436484
rect 504874 436450 504893 436484
rect 504821 436394 504893 436450
rect 504821 436360 504840 436394
rect 504874 436360 504893 436394
rect 504821 436304 504893 436360
rect 504821 436270 504840 436304
rect 504874 436270 504893 436304
rect 504821 436214 504893 436270
rect 504821 436180 504840 436214
rect 504874 436180 504893 436214
rect 505711 436866 505730 436900
rect 505764 436866 505783 436900
rect 505711 436810 505783 436866
rect 505711 436776 505730 436810
rect 505764 436776 505783 436810
rect 505711 436720 505783 436776
rect 505711 436686 505730 436720
rect 505764 436686 505783 436720
rect 505711 436630 505783 436686
rect 505711 436596 505730 436630
rect 505764 436596 505783 436630
rect 505711 436540 505783 436596
rect 505711 436506 505730 436540
rect 505764 436506 505783 436540
rect 505711 436450 505783 436506
rect 505711 436416 505730 436450
rect 505764 436416 505783 436450
rect 505711 436360 505783 436416
rect 505711 436326 505730 436360
rect 505764 436326 505783 436360
rect 505711 436270 505783 436326
rect 505711 436236 505730 436270
rect 505764 436236 505783 436270
rect 504821 436141 504893 436180
rect 505711 436180 505783 436236
rect 505711 436146 505730 436180
rect 505764 436146 505783 436180
rect 505711 436141 505783 436146
rect 504821 436122 505783 436141
rect 504821 436088 504934 436122
rect 504968 436088 505024 436122
rect 505058 436088 505114 436122
rect 505148 436088 505204 436122
rect 505238 436088 505294 436122
rect 505328 436088 505384 436122
rect 505418 436088 505474 436122
rect 505508 436088 505564 436122
rect 505598 436088 505654 436122
rect 505688 436088 505783 436122
rect 504821 436069 505783 436088
rect 506109 437012 507071 437031
rect 506109 436978 506241 437012
rect 506275 436978 506331 437012
rect 506365 436978 506421 437012
rect 506455 436978 506511 437012
rect 506545 436978 506601 437012
rect 506635 436978 506691 437012
rect 506725 436978 506781 437012
rect 506815 436978 506871 437012
rect 506905 436978 506961 437012
rect 506995 436978 507071 437012
rect 506109 436959 507071 436978
rect 506109 436934 506181 436959
rect 506109 436900 506128 436934
rect 506162 436900 506181 436934
rect 506109 436844 506181 436900
rect 506999 436900 507071 436959
rect 506109 436810 506128 436844
rect 506162 436810 506181 436844
rect 506109 436754 506181 436810
rect 506109 436720 506128 436754
rect 506162 436720 506181 436754
rect 506109 436664 506181 436720
rect 506109 436630 506128 436664
rect 506162 436630 506181 436664
rect 506109 436574 506181 436630
rect 506109 436540 506128 436574
rect 506162 436540 506181 436574
rect 506109 436484 506181 436540
rect 506109 436450 506128 436484
rect 506162 436450 506181 436484
rect 506109 436394 506181 436450
rect 506109 436360 506128 436394
rect 506162 436360 506181 436394
rect 506109 436304 506181 436360
rect 506109 436270 506128 436304
rect 506162 436270 506181 436304
rect 506109 436214 506181 436270
rect 506109 436180 506128 436214
rect 506162 436180 506181 436214
rect 506999 436866 507018 436900
rect 507052 436866 507071 436900
rect 506999 436810 507071 436866
rect 506999 436776 507018 436810
rect 507052 436776 507071 436810
rect 506999 436720 507071 436776
rect 506999 436686 507018 436720
rect 507052 436686 507071 436720
rect 506999 436630 507071 436686
rect 506999 436596 507018 436630
rect 507052 436596 507071 436630
rect 506999 436540 507071 436596
rect 506999 436506 507018 436540
rect 507052 436506 507071 436540
rect 506999 436450 507071 436506
rect 506999 436416 507018 436450
rect 507052 436416 507071 436450
rect 506999 436360 507071 436416
rect 506999 436326 507018 436360
rect 507052 436326 507071 436360
rect 506999 436270 507071 436326
rect 506999 436236 507018 436270
rect 507052 436236 507071 436270
rect 506109 436141 506181 436180
rect 506999 436180 507071 436236
rect 506999 436146 507018 436180
rect 507052 436146 507071 436180
rect 506999 436141 507071 436146
rect 506109 436122 507071 436141
rect 506109 436088 506222 436122
rect 506256 436088 506312 436122
rect 506346 436088 506402 436122
rect 506436 436088 506492 436122
rect 506526 436088 506582 436122
rect 506616 436088 506672 436122
rect 506706 436088 506762 436122
rect 506796 436088 506852 436122
rect 506886 436088 506942 436122
rect 506976 436088 507071 436122
rect 506109 436069 507071 436088
rect 507397 437012 508359 437031
rect 507397 436978 507529 437012
rect 507563 436978 507619 437012
rect 507653 436978 507709 437012
rect 507743 436978 507799 437012
rect 507833 436978 507889 437012
rect 507923 436978 507979 437012
rect 508013 436978 508069 437012
rect 508103 436978 508159 437012
rect 508193 436978 508249 437012
rect 508283 436978 508359 437012
rect 507397 436959 508359 436978
rect 507397 436934 507469 436959
rect 507397 436900 507416 436934
rect 507450 436900 507469 436934
rect 507397 436844 507469 436900
rect 508287 436900 508359 436959
rect 507397 436810 507416 436844
rect 507450 436810 507469 436844
rect 507397 436754 507469 436810
rect 507397 436720 507416 436754
rect 507450 436720 507469 436754
rect 507397 436664 507469 436720
rect 507397 436630 507416 436664
rect 507450 436630 507469 436664
rect 507397 436574 507469 436630
rect 507397 436540 507416 436574
rect 507450 436540 507469 436574
rect 507397 436484 507469 436540
rect 507397 436450 507416 436484
rect 507450 436450 507469 436484
rect 507397 436394 507469 436450
rect 507397 436360 507416 436394
rect 507450 436360 507469 436394
rect 507397 436304 507469 436360
rect 507397 436270 507416 436304
rect 507450 436270 507469 436304
rect 507397 436214 507469 436270
rect 507397 436180 507416 436214
rect 507450 436180 507469 436214
rect 508287 436866 508306 436900
rect 508340 436866 508359 436900
rect 508287 436810 508359 436866
rect 508287 436776 508306 436810
rect 508340 436776 508359 436810
rect 508287 436720 508359 436776
rect 508287 436686 508306 436720
rect 508340 436686 508359 436720
rect 508287 436630 508359 436686
rect 508287 436596 508306 436630
rect 508340 436596 508359 436630
rect 508287 436540 508359 436596
rect 508287 436506 508306 436540
rect 508340 436506 508359 436540
rect 508287 436450 508359 436506
rect 508287 436416 508306 436450
rect 508340 436416 508359 436450
rect 508287 436360 508359 436416
rect 508287 436326 508306 436360
rect 508340 436326 508359 436360
rect 508287 436270 508359 436326
rect 508287 436236 508306 436270
rect 508340 436236 508359 436270
rect 507397 436141 507469 436180
rect 508287 436180 508359 436236
rect 508287 436146 508306 436180
rect 508340 436146 508359 436180
rect 508287 436141 508359 436146
rect 507397 436122 508359 436141
rect 507397 436088 507510 436122
rect 507544 436088 507600 436122
rect 507634 436088 507690 436122
rect 507724 436088 507780 436122
rect 507814 436088 507870 436122
rect 507904 436088 507960 436122
rect 507994 436088 508050 436122
rect 508084 436088 508140 436122
rect 508174 436088 508230 436122
rect 508264 436088 508359 436122
rect 507397 436069 508359 436088
rect 508685 437012 509647 437031
rect 508685 436978 508817 437012
rect 508851 436978 508907 437012
rect 508941 436978 508997 437012
rect 509031 436978 509087 437012
rect 509121 436978 509177 437012
rect 509211 436978 509267 437012
rect 509301 436978 509357 437012
rect 509391 436978 509447 437012
rect 509481 436978 509537 437012
rect 509571 436978 509647 437012
rect 508685 436959 509647 436978
rect 508685 436934 508757 436959
rect 508685 436900 508704 436934
rect 508738 436900 508757 436934
rect 508685 436844 508757 436900
rect 509575 436900 509647 436959
rect 508685 436810 508704 436844
rect 508738 436810 508757 436844
rect 508685 436754 508757 436810
rect 508685 436720 508704 436754
rect 508738 436720 508757 436754
rect 508685 436664 508757 436720
rect 508685 436630 508704 436664
rect 508738 436630 508757 436664
rect 508685 436574 508757 436630
rect 508685 436540 508704 436574
rect 508738 436540 508757 436574
rect 508685 436484 508757 436540
rect 508685 436450 508704 436484
rect 508738 436450 508757 436484
rect 508685 436394 508757 436450
rect 508685 436360 508704 436394
rect 508738 436360 508757 436394
rect 508685 436304 508757 436360
rect 508685 436270 508704 436304
rect 508738 436270 508757 436304
rect 508685 436214 508757 436270
rect 508685 436180 508704 436214
rect 508738 436180 508757 436214
rect 509575 436866 509594 436900
rect 509628 436866 509647 436900
rect 509575 436810 509647 436866
rect 509575 436776 509594 436810
rect 509628 436776 509647 436810
rect 509575 436720 509647 436776
rect 509575 436686 509594 436720
rect 509628 436686 509647 436720
rect 509575 436630 509647 436686
rect 509575 436596 509594 436630
rect 509628 436596 509647 436630
rect 509575 436540 509647 436596
rect 509575 436506 509594 436540
rect 509628 436506 509647 436540
rect 509575 436450 509647 436506
rect 509575 436416 509594 436450
rect 509628 436416 509647 436450
rect 509575 436360 509647 436416
rect 509575 436326 509594 436360
rect 509628 436326 509647 436360
rect 509575 436270 509647 436326
rect 509575 436236 509594 436270
rect 509628 436236 509647 436270
rect 508685 436141 508757 436180
rect 509575 436180 509647 436236
rect 509575 436146 509594 436180
rect 509628 436146 509647 436180
rect 509575 436141 509647 436146
rect 508685 436122 509647 436141
rect 508685 436088 508798 436122
rect 508832 436088 508888 436122
rect 508922 436088 508978 436122
rect 509012 436088 509068 436122
rect 509102 436088 509158 436122
rect 509192 436088 509248 436122
rect 509282 436088 509338 436122
rect 509372 436088 509428 436122
rect 509462 436088 509518 436122
rect 509552 436088 509647 436122
rect 508685 436069 509647 436088
rect 509973 437012 510935 437031
rect 509973 436978 510105 437012
rect 510139 436978 510195 437012
rect 510229 436978 510285 437012
rect 510319 436978 510375 437012
rect 510409 436978 510465 437012
rect 510499 436978 510555 437012
rect 510589 436978 510645 437012
rect 510679 436978 510735 437012
rect 510769 436978 510825 437012
rect 510859 436978 510935 437012
rect 509973 436959 510935 436978
rect 509973 436934 510045 436959
rect 509973 436900 509992 436934
rect 510026 436900 510045 436934
rect 509973 436844 510045 436900
rect 510863 436900 510935 436959
rect 509973 436810 509992 436844
rect 510026 436810 510045 436844
rect 509973 436754 510045 436810
rect 509973 436720 509992 436754
rect 510026 436720 510045 436754
rect 509973 436664 510045 436720
rect 509973 436630 509992 436664
rect 510026 436630 510045 436664
rect 509973 436574 510045 436630
rect 509973 436540 509992 436574
rect 510026 436540 510045 436574
rect 509973 436484 510045 436540
rect 509973 436450 509992 436484
rect 510026 436450 510045 436484
rect 509973 436394 510045 436450
rect 509973 436360 509992 436394
rect 510026 436360 510045 436394
rect 509973 436304 510045 436360
rect 509973 436270 509992 436304
rect 510026 436270 510045 436304
rect 509973 436214 510045 436270
rect 509973 436180 509992 436214
rect 510026 436180 510045 436214
rect 510863 436866 510882 436900
rect 510916 436866 510935 436900
rect 510863 436810 510935 436866
rect 510863 436776 510882 436810
rect 510916 436776 510935 436810
rect 510863 436720 510935 436776
rect 510863 436686 510882 436720
rect 510916 436686 510935 436720
rect 510863 436630 510935 436686
rect 510863 436596 510882 436630
rect 510916 436596 510935 436630
rect 510863 436540 510935 436596
rect 510863 436506 510882 436540
rect 510916 436506 510935 436540
rect 510863 436450 510935 436506
rect 510863 436416 510882 436450
rect 510916 436416 510935 436450
rect 510863 436360 510935 436416
rect 510863 436326 510882 436360
rect 510916 436326 510935 436360
rect 510863 436270 510935 436326
rect 510863 436236 510882 436270
rect 510916 436236 510935 436270
rect 509973 436141 510045 436180
rect 510863 436180 510935 436236
rect 510863 436146 510882 436180
rect 510916 436146 510935 436180
rect 510863 436141 510935 436146
rect 509973 436122 510935 436141
rect 509973 436088 510086 436122
rect 510120 436088 510176 436122
rect 510210 436088 510266 436122
rect 510300 436088 510356 436122
rect 510390 436088 510446 436122
rect 510480 436088 510536 436122
rect 510570 436088 510626 436122
rect 510660 436088 510716 436122
rect 510750 436088 510806 436122
rect 510840 436088 510935 436122
rect 509973 436069 510935 436088
rect 511261 437012 512223 437031
rect 511261 436978 511393 437012
rect 511427 436978 511483 437012
rect 511517 436978 511573 437012
rect 511607 436978 511663 437012
rect 511697 436978 511753 437012
rect 511787 436978 511843 437012
rect 511877 436978 511933 437012
rect 511967 436978 512023 437012
rect 512057 436978 512113 437012
rect 512147 436978 512223 437012
rect 511261 436959 512223 436978
rect 511261 436934 511333 436959
rect 511261 436900 511280 436934
rect 511314 436900 511333 436934
rect 511261 436844 511333 436900
rect 512151 436900 512223 436959
rect 511261 436810 511280 436844
rect 511314 436810 511333 436844
rect 511261 436754 511333 436810
rect 511261 436720 511280 436754
rect 511314 436720 511333 436754
rect 511261 436664 511333 436720
rect 511261 436630 511280 436664
rect 511314 436630 511333 436664
rect 511261 436574 511333 436630
rect 511261 436540 511280 436574
rect 511314 436540 511333 436574
rect 511261 436484 511333 436540
rect 511261 436450 511280 436484
rect 511314 436450 511333 436484
rect 511261 436394 511333 436450
rect 511261 436360 511280 436394
rect 511314 436360 511333 436394
rect 511261 436304 511333 436360
rect 511261 436270 511280 436304
rect 511314 436270 511333 436304
rect 511261 436214 511333 436270
rect 511261 436180 511280 436214
rect 511314 436180 511333 436214
rect 512151 436866 512170 436900
rect 512204 436866 512223 436900
rect 512151 436810 512223 436866
rect 512151 436776 512170 436810
rect 512204 436776 512223 436810
rect 512151 436720 512223 436776
rect 512151 436686 512170 436720
rect 512204 436686 512223 436720
rect 512151 436630 512223 436686
rect 512151 436596 512170 436630
rect 512204 436596 512223 436630
rect 512151 436540 512223 436596
rect 512151 436506 512170 436540
rect 512204 436506 512223 436540
rect 512151 436450 512223 436506
rect 512151 436416 512170 436450
rect 512204 436416 512223 436450
rect 512151 436360 512223 436416
rect 512151 436326 512170 436360
rect 512204 436326 512223 436360
rect 512151 436270 512223 436326
rect 512151 436236 512170 436270
rect 512204 436236 512223 436270
rect 511261 436141 511333 436180
rect 512151 436180 512223 436236
rect 512151 436146 512170 436180
rect 512204 436146 512223 436180
rect 512151 436141 512223 436146
rect 511261 436122 512223 436141
rect 511261 436088 511374 436122
rect 511408 436088 511464 436122
rect 511498 436088 511554 436122
rect 511588 436088 511644 436122
rect 511678 436088 511734 436122
rect 511768 436088 511824 436122
rect 511858 436088 511914 436122
rect 511948 436088 512004 436122
rect 512038 436088 512094 436122
rect 512128 436088 512223 436122
rect 511261 436069 512223 436088
rect 512549 437012 513511 437031
rect 512549 436978 512681 437012
rect 512715 436978 512771 437012
rect 512805 436978 512861 437012
rect 512895 436978 512951 437012
rect 512985 436978 513041 437012
rect 513075 436978 513131 437012
rect 513165 436978 513221 437012
rect 513255 436978 513311 437012
rect 513345 436978 513401 437012
rect 513435 436978 513511 437012
rect 512549 436959 513511 436978
rect 512549 436934 512621 436959
rect 512549 436900 512568 436934
rect 512602 436900 512621 436934
rect 512549 436844 512621 436900
rect 513439 436900 513511 436959
rect 512549 436810 512568 436844
rect 512602 436810 512621 436844
rect 512549 436754 512621 436810
rect 512549 436720 512568 436754
rect 512602 436720 512621 436754
rect 512549 436664 512621 436720
rect 512549 436630 512568 436664
rect 512602 436630 512621 436664
rect 512549 436574 512621 436630
rect 512549 436540 512568 436574
rect 512602 436540 512621 436574
rect 512549 436484 512621 436540
rect 512549 436450 512568 436484
rect 512602 436450 512621 436484
rect 512549 436394 512621 436450
rect 512549 436360 512568 436394
rect 512602 436360 512621 436394
rect 512549 436304 512621 436360
rect 512549 436270 512568 436304
rect 512602 436270 512621 436304
rect 512549 436214 512621 436270
rect 512549 436180 512568 436214
rect 512602 436180 512621 436214
rect 513439 436866 513458 436900
rect 513492 436866 513511 436900
rect 513439 436810 513511 436866
rect 513439 436776 513458 436810
rect 513492 436776 513511 436810
rect 513439 436720 513511 436776
rect 513439 436686 513458 436720
rect 513492 436686 513511 436720
rect 513439 436630 513511 436686
rect 513439 436596 513458 436630
rect 513492 436596 513511 436630
rect 513439 436540 513511 436596
rect 513439 436506 513458 436540
rect 513492 436506 513511 436540
rect 513439 436450 513511 436506
rect 513439 436416 513458 436450
rect 513492 436416 513511 436450
rect 513439 436360 513511 436416
rect 513439 436326 513458 436360
rect 513492 436326 513511 436360
rect 513439 436270 513511 436326
rect 513439 436236 513458 436270
rect 513492 436236 513511 436270
rect 512549 436141 512621 436180
rect 513439 436180 513511 436236
rect 513439 436146 513458 436180
rect 513492 436146 513511 436180
rect 513439 436141 513511 436146
rect 512549 436122 513511 436141
rect 512549 436088 512662 436122
rect 512696 436088 512752 436122
rect 512786 436088 512842 436122
rect 512876 436088 512932 436122
rect 512966 436088 513022 436122
rect 513056 436088 513112 436122
rect 513146 436088 513202 436122
rect 513236 436088 513292 436122
rect 513326 436088 513382 436122
rect 513416 436088 513511 436122
rect 512549 436069 513511 436088
rect 503533 435724 504495 435743
rect 503533 435690 503665 435724
rect 503699 435690 503755 435724
rect 503789 435690 503845 435724
rect 503879 435690 503935 435724
rect 503969 435690 504025 435724
rect 504059 435690 504115 435724
rect 504149 435690 504205 435724
rect 504239 435690 504295 435724
rect 504329 435690 504385 435724
rect 504419 435690 504495 435724
rect 503533 435671 504495 435690
rect 503533 435646 503605 435671
rect 503533 435612 503552 435646
rect 503586 435612 503605 435646
rect 503533 435556 503605 435612
rect 504423 435612 504495 435671
rect 503533 435522 503552 435556
rect 503586 435522 503605 435556
rect 503533 435466 503605 435522
rect 503533 435432 503552 435466
rect 503586 435432 503605 435466
rect 503533 435376 503605 435432
rect 503533 435342 503552 435376
rect 503586 435342 503605 435376
rect 503533 435286 503605 435342
rect 503533 435252 503552 435286
rect 503586 435252 503605 435286
rect 503533 435196 503605 435252
rect 503533 435162 503552 435196
rect 503586 435162 503605 435196
rect 503533 435106 503605 435162
rect 503533 435072 503552 435106
rect 503586 435072 503605 435106
rect 503533 435016 503605 435072
rect 503533 434982 503552 435016
rect 503586 434982 503605 435016
rect 503533 434926 503605 434982
rect 503533 434892 503552 434926
rect 503586 434892 503605 434926
rect 504423 435578 504442 435612
rect 504476 435578 504495 435612
rect 504423 435522 504495 435578
rect 504423 435488 504442 435522
rect 504476 435488 504495 435522
rect 504423 435432 504495 435488
rect 504423 435398 504442 435432
rect 504476 435398 504495 435432
rect 504423 435342 504495 435398
rect 504423 435308 504442 435342
rect 504476 435308 504495 435342
rect 504423 435252 504495 435308
rect 504423 435218 504442 435252
rect 504476 435218 504495 435252
rect 504423 435162 504495 435218
rect 504423 435128 504442 435162
rect 504476 435128 504495 435162
rect 504423 435072 504495 435128
rect 504423 435038 504442 435072
rect 504476 435038 504495 435072
rect 504423 434982 504495 435038
rect 504423 434948 504442 434982
rect 504476 434948 504495 434982
rect 503533 434853 503605 434892
rect 504423 434892 504495 434948
rect 504423 434858 504442 434892
rect 504476 434858 504495 434892
rect 504423 434853 504495 434858
rect 503533 434834 504495 434853
rect 503533 434800 503646 434834
rect 503680 434800 503736 434834
rect 503770 434800 503826 434834
rect 503860 434800 503916 434834
rect 503950 434800 504006 434834
rect 504040 434800 504096 434834
rect 504130 434800 504186 434834
rect 504220 434800 504276 434834
rect 504310 434800 504366 434834
rect 504400 434800 504495 434834
rect 503533 434781 504495 434800
rect 504821 435724 505783 435743
rect 504821 435690 504953 435724
rect 504987 435690 505043 435724
rect 505077 435690 505133 435724
rect 505167 435690 505223 435724
rect 505257 435690 505313 435724
rect 505347 435690 505403 435724
rect 505437 435690 505493 435724
rect 505527 435690 505583 435724
rect 505617 435690 505673 435724
rect 505707 435690 505783 435724
rect 504821 435671 505783 435690
rect 504821 435646 504893 435671
rect 504821 435612 504840 435646
rect 504874 435612 504893 435646
rect 504821 435556 504893 435612
rect 505711 435612 505783 435671
rect 504821 435522 504840 435556
rect 504874 435522 504893 435556
rect 504821 435466 504893 435522
rect 504821 435432 504840 435466
rect 504874 435432 504893 435466
rect 504821 435376 504893 435432
rect 504821 435342 504840 435376
rect 504874 435342 504893 435376
rect 504821 435286 504893 435342
rect 504821 435252 504840 435286
rect 504874 435252 504893 435286
rect 504821 435196 504893 435252
rect 504821 435162 504840 435196
rect 504874 435162 504893 435196
rect 504821 435106 504893 435162
rect 504821 435072 504840 435106
rect 504874 435072 504893 435106
rect 504821 435016 504893 435072
rect 504821 434982 504840 435016
rect 504874 434982 504893 435016
rect 504821 434926 504893 434982
rect 504821 434892 504840 434926
rect 504874 434892 504893 434926
rect 505711 435578 505730 435612
rect 505764 435578 505783 435612
rect 505711 435522 505783 435578
rect 505711 435488 505730 435522
rect 505764 435488 505783 435522
rect 505711 435432 505783 435488
rect 505711 435398 505730 435432
rect 505764 435398 505783 435432
rect 505711 435342 505783 435398
rect 505711 435308 505730 435342
rect 505764 435308 505783 435342
rect 505711 435252 505783 435308
rect 505711 435218 505730 435252
rect 505764 435218 505783 435252
rect 505711 435162 505783 435218
rect 505711 435128 505730 435162
rect 505764 435128 505783 435162
rect 505711 435072 505783 435128
rect 505711 435038 505730 435072
rect 505764 435038 505783 435072
rect 505711 434982 505783 435038
rect 505711 434948 505730 434982
rect 505764 434948 505783 434982
rect 504821 434853 504893 434892
rect 505711 434892 505783 434948
rect 505711 434858 505730 434892
rect 505764 434858 505783 434892
rect 505711 434853 505783 434858
rect 504821 434834 505783 434853
rect 504821 434800 504934 434834
rect 504968 434800 505024 434834
rect 505058 434800 505114 434834
rect 505148 434800 505204 434834
rect 505238 434800 505294 434834
rect 505328 434800 505384 434834
rect 505418 434800 505474 434834
rect 505508 434800 505564 434834
rect 505598 434800 505654 434834
rect 505688 434800 505783 434834
rect 504821 434781 505783 434800
rect 506109 435724 507071 435743
rect 506109 435690 506241 435724
rect 506275 435690 506331 435724
rect 506365 435690 506421 435724
rect 506455 435690 506511 435724
rect 506545 435690 506601 435724
rect 506635 435690 506691 435724
rect 506725 435690 506781 435724
rect 506815 435690 506871 435724
rect 506905 435690 506961 435724
rect 506995 435690 507071 435724
rect 506109 435671 507071 435690
rect 506109 435646 506181 435671
rect 506109 435612 506128 435646
rect 506162 435612 506181 435646
rect 506109 435556 506181 435612
rect 506999 435612 507071 435671
rect 506109 435522 506128 435556
rect 506162 435522 506181 435556
rect 506109 435466 506181 435522
rect 506109 435432 506128 435466
rect 506162 435432 506181 435466
rect 506109 435376 506181 435432
rect 506109 435342 506128 435376
rect 506162 435342 506181 435376
rect 506109 435286 506181 435342
rect 506109 435252 506128 435286
rect 506162 435252 506181 435286
rect 506109 435196 506181 435252
rect 506109 435162 506128 435196
rect 506162 435162 506181 435196
rect 506109 435106 506181 435162
rect 506109 435072 506128 435106
rect 506162 435072 506181 435106
rect 506109 435016 506181 435072
rect 506109 434982 506128 435016
rect 506162 434982 506181 435016
rect 506109 434926 506181 434982
rect 506109 434892 506128 434926
rect 506162 434892 506181 434926
rect 506999 435578 507018 435612
rect 507052 435578 507071 435612
rect 506999 435522 507071 435578
rect 506999 435488 507018 435522
rect 507052 435488 507071 435522
rect 506999 435432 507071 435488
rect 506999 435398 507018 435432
rect 507052 435398 507071 435432
rect 506999 435342 507071 435398
rect 506999 435308 507018 435342
rect 507052 435308 507071 435342
rect 506999 435252 507071 435308
rect 506999 435218 507018 435252
rect 507052 435218 507071 435252
rect 506999 435162 507071 435218
rect 506999 435128 507018 435162
rect 507052 435128 507071 435162
rect 506999 435072 507071 435128
rect 506999 435038 507018 435072
rect 507052 435038 507071 435072
rect 506999 434982 507071 435038
rect 506999 434948 507018 434982
rect 507052 434948 507071 434982
rect 506109 434853 506181 434892
rect 506999 434892 507071 434948
rect 506999 434858 507018 434892
rect 507052 434858 507071 434892
rect 506999 434853 507071 434858
rect 506109 434834 507071 434853
rect 506109 434800 506222 434834
rect 506256 434800 506312 434834
rect 506346 434800 506402 434834
rect 506436 434800 506492 434834
rect 506526 434800 506582 434834
rect 506616 434800 506672 434834
rect 506706 434800 506762 434834
rect 506796 434800 506852 434834
rect 506886 434800 506942 434834
rect 506976 434800 507071 434834
rect 506109 434781 507071 434800
rect 507397 435724 508359 435743
rect 507397 435690 507529 435724
rect 507563 435690 507619 435724
rect 507653 435690 507709 435724
rect 507743 435690 507799 435724
rect 507833 435690 507889 435724
rect 507923 435690 507979 435724
rect 508013 435690 508069 435724
rect 508103 435690 508159 435724
rect 508193 435690 508249 435724
rect 508283 435690 508359 435724
rect 507397 435671 508359 435690
rect 507397 435646 507469 435671
rect 507397 435612 507416 435646
rect 507450 435612 507469 435646
rect 507397 435556 507469 435612
rect 508287 435612 508359 435671
rect 507397 435522 507416 435556
rect 507450 435522 507469 435556
rect 507397 435466 507469 435522
rect 507397 435432 507416 435466
rect 507450 435432 507469 435466
rect 507397 435376 507469 435432
rect 507397 435342 507416 435376
rect 507450 435342 507469 435376
rect 507397 435286 507469 435342
rect 507397 435252 507416 435286
rect 507450 435252 507469 435286
rect 507397 435196 507469 435252
rect 507397 435162 507416 435196
rect 507450 435162 507469 435196
rect 507397 435106 507469 435162
rect 507397 435072 507416 435106
rect 507450 435072 507469 435106
rect 507397 435016 507469 435072
rect 507397 434982 507416 435016
rect 507450 434982 507469 435016
rect 507397 434926 507469 434982
rect 507397 434892 507416 434926
rect 507450 434892 507469 434926
rect 508287 435578 508306 435612
rect 508340 435578 508359 435612
rect 508287 435522 508359 435578
rect 508287 435488 508306 435522
rect 508340 435488 508359 435522
rect 508287 435432 508359 435488
rect 508287 435398 508306 435432
rect 508340 435398 508359 435432
rect 508287 435342 508359 435398
rect 508287 435308 508306 435342
rect 508340 435308 508359 435342
rect 508287 435252 508359 435308
rect 508287 435218 508306 435252
rect 508340 435218 508359 435252
rect 508287 435162 508359 435218
rect 508287 435128 508306 435162
rect 508340 435128 508359 435162
rect 508287 435072 508359 435128
rect 508287 435038 508306 435072
rect 508340 435038 508359 435072
rect 508287 434982 508359 435038
rect 508287 434948 508306 434982
rect 508340 434948 508359 434982
rect 507397 434853 507469 434892
rect 508287 434892 508359 434948
rect 508287 434858 508306 434892
rect 508340 434858 508359 434892
rect 508287 434853 508359 434858
rect 507397 434834 508359 434853
rect 507397 434800 507510 434834
rect 507544 434800 507600 434834
rect 507634 434800 507690 434834
rect 507724 434800 507780 434834
rect 507814 434800 507870 434834
rect 507904 434800 507960 434834
rect 507994 434800 508050 434834
rect 508084 434800 508140 434834
rect 508174 434800 508230 434834
rect 508264 434800 508359 434834
rect 507397 434781 508359 434800
rect 508685 435724 509647 435743
rect 508685 435690 508817 435724
rect 508851 435690 508907 435724
rect 508941 435690 508997 435724
rect 509031 435690 509087 435724
rect 509121 435690 509177 435724
rect 509211 435690 509267 435724
rect 509301 435690 509357 435724
rect 509391 435690 509447 435724
rect 509481 435690 509537 435724
rect 509571 435690 509647 435724
rect 508685 435671 509647 435690
rect 508685 435646 508757 435671
rect 508685 435612 508704 435646
rect 508738 435612 508757 435646
rect 508685 435556 508757 435612
rect 509575 435612 509647 435671
rect 508685 435522 508704 435556
rect 508738 435522 508757 435556
rect 508685 435466 508757 435522
rect 508685 435432 508704 435466
rect 508738 435432 508757 435466
rect 508685 435376 508757 435432
rect 508685 435342 508704 435376
rect 508738 435342 508757 435376
rect 508685 435286 508757 435342
rect 508685 435252 508704 435286
rect 508738 435252 508757 435286
rect 508685 435196 508757 435252
rect 508685 435162 508704 435196
rect 508738 435162 508757 435196
rect 508685 435106 508757 435162
rect 508685 435072 508704 435106
rect 508738 435072 508757 435106
rect 508685 435016 508757 435072
rect 508685 434982 508704 435016
rect 508738 434982 508757 435016
rect 508685 434926 508757 434982
rect 508685 434892 508704 434926
rect 508738 434892 508757 434926
rect 509575 435578 509594 435612
rect 509628 435578 509647 435612
rect 509575 435522 509647 435578
rect 509575 435488 509594 435522
rect 509628 435488 509647 435522
rect 509575 435432 509647 435488
rect 509575 435398 509594 435432
rect 509628 435398 509647 435432
rect 509575 435342 509647 435398
rect 509575 435308 509594 435342
rect 509628 435308 509647 435342
rect 509575 435252 509647 435308
rect 509575 435218 509594 435252
rect 509628 435218 509647 435252
rect 509575 435162 509647 435218
rect 509575 435128 509594 435162
rect 509628 435128 509647 435162
rect 509575 435072 509647 435128
rect 509575 435038 509594 435072
rect 509628 435038 509647 435072
rect 509575 434982 509647 435038
rect 509575 434948 509594 434982
rect 509628 434948 509647 434982
rect 508685 434853 508757 434892
rect 509575 434892 509647 434948
rect 509575 434858 509594 434892
rect 509628 434858 509647 434892
rect 509575 434853 509647 434858
rect 508685 434834 509647 434853
rect 508685 434800 508798 434834
rect 508832 434800 508888 434834
rect 508922 434800 508978 434834
rect 509012 434800 509068 434834
rect 509102 434800 509158 434834
rect 509192 434800 509248 434834
rect 509282 434800 509338 434834
rect 509372 434800 509428 434834
rect 509462 434800 509518 434834
rect 509552 434800 509647 434834
rect 508685 434781 509647 434800
rect 509973 435724 510935 435743
rect 509973 435690 510105 435724
rect 510139 435690 510195 435724
rect 510229 435690 510285 435724
rect 510319 435690 510375 435724
rect 510409 435690 510465 435724
rect 510499 435690 510555 435724
rect 510589 435690 510645 435724
rect 510679 435690 510735 435724
rect 510769 435690 510825 435724
rect 510859 435690 510935 435724
rect 509973 435671 510935 435690
rect 509973 435646 510045 435671
rect 509973 435612 509992 435646
rect 510026 435612 510045 435646
rect 509973 435556 510045 435612
rect 510863 435612 510935 435671
rect 509973 435522 509992 435556
rect 510026 435522 510045 435556
rect 509973 435466 510045 435522
rect 509973 435432 509992 435466
rect 510026 435432 510045 435466
rect 509973 435376 510045 435432
rect 509973 435342 509992 435376
rect 510026 435342 510045 435376
rect 509973 435286 510045 435342
rect 509973 435252 509992 435286
rect 510026 435252 510045 435286
rect 509973 435196 510045 435252
rect 509973 435162 509992 435196
rect 510026 435162 510045 435196
rect 509973 435106 510045 435162
rect 509973 435072 509992 435106
rect 510026 435072 510045 435106
rect 509973 435016 510045 435072
rect 509973 434982 509992 435016
rect 510026 434982 510045 435016
rect 509973 434926 510045 434982
rect 509973 434892 509992 434926
rect 510026 434892 510045 434926
rect 510863 435578 510882 435612
rect 510916 435578 510935 435612
rect 510863 435522 510935 435578
rect 510863 435488 510882 435522
rect 510916 435488 510935 435522
rect 510863 435432 510935 435488
rect 510863 435398 510882 435432
rect 510916 435398 510935 435432
rect 510863 435342 510935 435398
rect 510863 435308 510882 435342
rect 510916 435308 510935 435342
rect 510863 435252 510935 435308
rect 510863 435218 510882 435252
rect 510916 435218 510935 435252
rect 510863 435162 510935 435218
rect 510863 435128 510882 435162
rect 510916 435128 510935 435162
rect 510863 435072 510935 435128
rect 510863 435038 510882 435072
rect 510916 435038 510935 435072
rect 510863 434982 510935 435038
rect 510863 434948 510882 434982
rect 510916 434948 510935 434982
rect 509973 434853 510045 434892
rect 510863 434892 510935 434948
rect 510863 434858 510882 434892
rect 510916 434858 510935 434892
rect 510863 434853 510935 434858
rect 509973 434834 510935 434853
rect 509973 434800 510086 434834
rect 510120 434800 510176 434834
rect 510210 434800 510266 434834
rect 510300 434800 510356 434834
rect 510390 434800 510446 434834
rect 510480 434800 510536 434834
rect 510570 434800 510626 434834
rect 510660 434800 510716 434834
rect 510750 434800 510806 434834
rect 510840 434800 510935 434834
rect 509973 434781 510935 434800
rect 511261 435724 512223 435743
rect 511261 435690 511393 435724
rect 511427 435690 511483 435724
rect 511517 435690 511573 435724
rect 511607 435690 511663 435724
rect 511697 435690 511753 435724
rect 511787 435690 511843 435724
rect 511877 435690 511933 435724
rect 511967 435690 512023 435724
rect 512057 435690 512113 435724
rect 512147 435690 512223 435724
rect 511261 435671 512223 435690
rect 511261 435646 511333 435671
rect 511261 435612 511280 435646
rect 511314 435612 511333 435646
rect 511261 435556 511333 435612
rect 512151 435612 512223 435671
rect 511261 435522 511280 435556
rect 511314 435522 511333 435556
rect 511261 435466 511333 435522
rect 511261 435432 511280 435466
rect 511314 435432 511333 435466
rect 511261 435376 511333 435432
rect 511261 435342 511280 435376
rect 511314 435342 511333 435376
rect 511261 435286 511333 435342
rect 511261 435252 511280 435286
rect 511314 435252 511333 435286
rect 511261 435196 511333 435252
rect 511261 435162 511280 435196
rect 511314 435162 511333 435196
rect 511261 435106 511333 435162
rect 511261 435072 511280 435106
rect 511314 435072 511333 435106
rect 511261 435016 511333 435072
rect 511261 434982 511280 435016
rect 511314 434982 511333 435016
rect 511261 434926 511333 434982
rect 511261 434892 511280 434926
rect 511314 434892 511333 434926
rect 512151 435578 512170 435612
rect 512204 435578 512223 435612
rect 512151 435522 512223 435578
rect 512151 435488 512170 435522
rect 512204 435488 512223 435522
rect 512151 435432 512223 435488
rect 512151 435398 512170 435432
rect 512204 435398 512223 435432
rect 512151 435342 512223 435398
rect 512151 435308 512170 435342
rect 512204 435308 512223 435342
rect 512151 435252 512223 435308
rect 512151 435218 512170 435252
rect 512204 435218 512223 435252
rect 512151 435162 512223 435218
rect 512151 435128 512170 435162
rect 512204 435128 512223 435162
rect 512151 435072 512223 435128
rect 512151 435038 512170 435072
rect 512204 435038 512223 435072
rect 512151 434982 512223 435038
rect 512151 434948 512170 434982
rect 512204 434948 512223 434982
rect 511261 434853 511333 434892
rect 512151 434892 512223 434948
rect 512151 434858 512170 434892
rect 512204 434858 512223 434892
rect 512151 434853 512223 434858
rect 511261 434834 512223 434853
rect 511261 434800 511374 434834
rect 511408 434800 511464 434834
rect 511498 434800 511554 434834
rect 511588 434800 511644 434834
rect 511678 434800 511734 434834
rect 511768 434800 511824 434834
rect 511858 434800 511914 434834
rect 511948 434800 512004 434834
rect 512038 434800 512094 434834
rect 512128 434800 512223 434834
rect 511261 434781 512223 434800
rect 512549 435724 513511 435743
rect 512549 435690 512681 435724
rect 512715 435690 512771 435724
rect 512805 435690 512861 435724
rect 512895 435690 512951 435724
rect 512985 435690 513041 435724
rect 513075 435690 513131 435724
rect 513165 435690 513221 435724
rect 513255 435690 513311 435724
rect 513345 435690 513401 435724
rect 513435 435690 513511 435724
rect 512549 435671 513511 435690
rect 512549 435646 512621 435671
rect 512549 435612 512568 435646
rect 512602 435612 512621 435646
rect 512549 435556 512621 435612
rect 513439 435612 513511 435671
rect 512549 435522 512568 435556
rect 512602 435522 512621 435556
rect 512549 435466 512621 435522
rect 512549 435432 512568 435466
rect 512602 435432 512621 435466
rect 512549 435376 512621 435432
rect 512549 435342 512568 435376
rect 512602 435342 512621 435376
rect 512549 435286 512621 435342
rect 512549 435252 512568 435286
rect 512602 435252 512621 435286
rect 512549 435196 512621 435252
rect 512549 435162 512568 435196
rect 512602 435162 512621 435196
rect 512549 435106 512621 435162
rect 512549 435072 512568 435106
rect 512602 435072 512621 435106
rect 512549 435016 512621 435072
rect 512549 434982 512568 435016
rect 512602 434982 512621 435016
rect 512549 434926 512621 434982
rect 512549 434892 512568 434926
rect 512602 434892 512621 434926
rect 513439 435578 513458 435612
rect 513492 435578 513511 435612
rect 513439 435522 513511 435578
rect 513439 435488 513458 435522
rect 513492 435488 513511 435522
rect 513439 435432 513511 435488
rect 513439 435398 513458 435432
rect 513492 435398 513511 435432
rect 513439 435342 513511 435398
rect 513439 435308 513458 435342
rect 513492 435308 513511 435342
rect 513439 435252 513511 435308
rect 513439 435218 513458 435252
rect 513492 435218 513511 435252
rect 513439 435162 513511 435218
rect 513439 435128 513458 435162
rect 513492 435128 513511 435162
rect 513439 435072 513511 435128
rect 513439 435038 513458 435072
rect 513492 435038 513511 435072
rect 513439 434982 513511 435038
rect 513439 434948 513458 434982
rect 513492 434948 513511 434982
rect 512549 434853 512621 434892
rect 513439 434892 513511 434948
rect 513439 434858 513458 434892
rect 513492 434858 513511 434892
rect 513439 434853 513511 434858
rect 512549 434834 513511 434853
rect 512549 434800 512662 434834
rect 512696 434800 512752 434834
rect 512786 434800 512842 434834
rect 512876 434800 512932 434834
rect 512966 434800 513022 434834
rect 513056 434800 513112 434834
rect 513146 434800 513202 434834
rect 513236 434800 513292 434834
rect 513326 434800 513382 434834
rect 513416 434800 513511 434834
rect 512549 434781 513511 434800
rect 503533 434436 504495 434455
rect 503533 434402 503665 434436
rect 503699 434402 503755 434436
rect 503789 434402 503845 434436
rect 503879 434402 503935 434436
rect 503969 434402 504025 434436
rect 504059 434402 504115 434436
rect 504149 434402 504205 434436
rect 504239 434402 504295 434436
rect 504329 434402 504385 434436
rect 504419 434402 504495 434436
rect 503533 434383 504495 434402
rect 503533 434358 503605 434383
rect 503533 434324 503552 434358
rect 503586 434324 503605 434358
rect 503533 434268 503605 434324
rect 504423 434324 504495 434383
rect 503533 434234 503552 434268
rect 503586 434234 503605 434268
rect 503533 434178 503605 434234
rect 503533 434144 503552 434178
rect 503586 434144 503605 434178
rect 503533 434088 503605 434144
rect 503533 434054 503552 434088
rect 503586 434054 503605 434088
rect 503533 433998 503605 434054
rect 503533 433964 503552 433998
rect 503586 433964 503605 433998
rect 503533 433908 503605 433964
rect 503533 433874 503552 433908
rect 503586 433874 503605 433908
rect 503533 433818 503605 433874
rect 503533 433784 503552 433818
rect 503586 433784 503605 433818
rect 503533 433728 503605 433784
rect 503533 433694 503552 433728
rect 503586 433694 503605 433728
rect 503533 433638 503605 433694
rect 503533 433604 503552 433638
rect 503586 433604 503605 433638
rect 504423 434290 504442 434324
rect 504476 434290 504495 434324
rect 504423 434234 504495 434290
rect 504423 434200 504442 434234
rect 504476 434200 504495 434234
rect 504423 434144 504495 434200
rect 504423 434110 504442 434144
rect 504476 434110 504495 434144
rect 504423 434054 504495 434110
rect 504423 434020 504442 434054
rect 504476 434020 504495 434054
rect 504423 433964 504495 434020
rect 504423 433930 504442 433964
rect 504476 433930 504495 433964
rect 504423 433874 504495 433930
rect 504423 433840 504442 433874
rect 504476 433840 504495 433874
rect 504423 433784 504495 433840
rect 504423 433750 504442 433784
rect 504476 433750 504495 433784
rect 504423 433694 504495 433750
rect 504423 433660 504442 433694
rect 504476 433660 504495 433694
rect 503533 433565 503605 433604
rect 504423 433604 504495 433660
rect 504423 433570 504442 433604
rect 504476 433570 504495 433604
rect 504423 433565 504495 433570
rect 503533 433546 504495 433565
rect 503533 433512 503646 433546
rect 503680 433512 503736 433546
rect 503770 433512 503826 433546
rect 503860 433512 503916 433546
rect 503950 433512 504006 433546
rect 504040 433512 504096 433546
rect 504130 433512 504186 433546
rect 504220 433512 504276 433546
rect 504310 433512 504366 433546
rect 504400 433512 504495 433546
rect 503533 433493 504495 433512
rect 504821 434436 505783 434455
rect 504821 434402 504953 434436
rect 504987 434402 505043 434436
rect 505077 434402 505133 434436
rect 505167 434402 505223 434436
rect 505257 434402 505313 434436
rect 505347 434402 505403 434436
rect 505437 434402 505493 434436
rect 505527 434402 505583 434436
rect 505617 434402 505673 434436
rect 505707 434402 505783 434436
rect 504821 434383 505783 434402
rect 504821 434358 504893 434383
rect 504821 434324 504840 434358
rect 504874 434324 504893 434358
rect 504821 434268 504893 434324
rect 505711 434324 505783 434383
rect 504821 434234 504840 434268
rect 504874 434234 504893 434268
rect 504821 434178 504893 434234
rect 504821 434144 504840 434178
rect 504874 434144 504893 434178
rect 504821 434088 504893 434144
rect 504821 434054 504840 434088
rect 504874 434054 504893 434088
rect 504821 433998 504893 434054
rect 504821 433964 504840 433998
rect 504874 433964 504893 433998
rect 504821 433908 504893 433964
rect 504821 433874 504840 433908
rect 504874 433874 504893 433908
rect 504821 433818 504893 433874
rect 504821 433784 504840 433818
rect 504874 433784 504893 433818
rect 504821 433728 504893 433784
rect 504821 433694 504840 433728
rect 504874 433694 504893 433728
rect 504821 433638 504893 433694
rect 504821 433604 504840 433638
rect 504874 433604 504893 433638
rect 505711 434290 505730 434324
rect 505764 434290 505783 434324
rect 505711 434234 505783 434290
rect 505711 434200 505730 434234
rect 505764 434200 505783 434234
rect 505711 434144 505783 434200
rect 505711 434110 505730 434144
rect 505764 434110 505783 434144
rect 505711 434054 505783 434110
rect 505711 434020 505730 434054
rect 505764 434020 505783 434054
rect 505711 433964 505783 434020
rect 505711 433930 505730 433964
rect 505764 433930 505783 433964
rect 505711 433874 505783 433930
rect 505711 433840 505730 433874
rect 505764 433840 505783 433874
rect 505711 433784 505783 433840
rect 505711 433750 505730 433784
rect 505764 433750 505783 433784
rect 505711 433694 505783 433750
rect 505711 433660 505730 433694
rect 505764 433660 505783 433694
rect 504821 433565 504893 433604
rect 505711 433604 505783 433660
rect 505711 433570 505730 433604
rect 505764 433570 505783 433604
rect 505711 433565 505783 433570
rect 504821 433546 505783 433565
rect 504821 433512 504934 433546
rect 504968 433512 505024 433546
rect 505058 433512 505114 433546
rect 505148 433512 505204 433546
rect 505238 433512 505294 433546
rect 505328 433512 505384 433546
rect 505418 433512 505474 433546
rect 505508 433512 505564 433546
rect 505598 433512 505654 433546
rect 505688 433512 505783 433546
rect 504821 433493 505783 433512
rect 506109 434436 507071 434455
rect 506109 434402 506241 434436
rect 506275 434402 506331 434436
rect 506365 434402 506421 434436
rect 506455 434402 506511 434436
rect 506545 434402 506601 434436
rect 506635 434402 506691 434436
rect 506725 434402 506781 434436
rect 506815 434402 506871 434436
rect 506905 434402 506961 434436
rect 506995 434402 507071 434436
rect 506109 434383 507071 434402
rect 506109 434358 506181 434383
rect 506109 434324 506128 434358
rect 506162 434324 506181 434358
rect 506109 434268 506181 434324
rect 506999 434324 507071 434383
rect 506109 434234 506128 434268
rect 506162 434234 506181 434268
rect 506109 434178 506181 434234
rect 506109 434144 506128 434178
rect 506162 434144 506181 434178
rect 506109 434088 506181 434144
rect 506109 434054 506128 434088
rect 506162 434054 506181 434088
rect 506109 433998 506181 434054
rect 506109 433964 506128 433998
rect 506162 433964 506181 433998
rect 506109 433908 506181 433964
rect 506109 433874 506128 433908
rect 506162 433874 506181 433908
rect 506109 433818 506181 433874
rect 506109 433784 506128 433818
rect 506162 433784 506181 433818
rect 506109 433728 506181 433784
rect 506109 433694 506128 433728
rect 506162 433694 506181 433728
rect 506109 433638 506181 433694
rect 506109 433604 506128 433638
rect 506162 433604 506181 433638
rect 506999 434290 507018 434324
rect 507052 434290 507071 434324
rect 506999 434234 507071 434290
rect 506999 434200 507018 434234
rect 507052 434200 507071 434234
rect 506999 434144 507071 434200
rect 506999 434110 507018 434144
rect 507052 434110 507071 434144
rect 506999 434054 507071 434110
rect 506999 434020 507018 434054
rect 507052 434020 507071 434054
rect 506999 433964 507071 434020
rect 506999 433930 507018 433964
rect 507052 433930 507071 433964
rect 506999 433874 507071 433930
rect 506999 433840 507018 433874
rect 507052 433840 507071 433874
rect 506999 433784 507071 433840
rect 506999 433750 507018 433784
rect 507052 433750 507071 433784
rect 506999 433694 507071 433750
rect 506999 433660 507018 433694
rect 507052 433660 507071 433694
rect 506109 433565 506181 433604
rect 506999 433604 507071 433660
rect 506999 433570 507018 433604
rect 507052 433570 507071 433604
rect 506999 433565 507071 433570
rect 506109 433546 507071 433565
rect 506109 433512 506222 433546
rect 506256 433512 506312 433546
rect 506346 433512 506402 433546
rect 506436 433512 506492 433546
rect 506526 433512 506582 433546
rect 506616 433512 506672 433546
rect 506706 433512 506762 433546
rect 506796 433512 506852 433546
rect 506886 433512 506942 433546
rect 506976 433512 507071 433546
rect 506109 433493 507071 433512
rect 507397 434436 508359 434455
rect 507397 434402 507529 434436
rect 507563 434402 507619 434436
rect 507653 434402 507709 434436
rect 507743 434402 507799 434436
rect 507833 434402 507889 434436
rect 507923 434402 507979 434436
rect 508013 434402 508069 434436
rect 508103 434402 508159 434436
rect 508193 434402 508249 434436
rect 508283 434402 508359 434436
rect 507397 434383 508359 434402
rect 507397 434358 507469 434383
rect 507397 434324 507416 434358
rect 507450 434324 507469 434358
rect 507397 434268 507469 434324
rect 508287 434324 508359 434383
rect 507397 434234 507416 434268
rect 507450 434234 507469 434268
rect 507397 434178 507469 434234
rect 507397 434144 507416 434178
rect 507450 434144 507469 434178
rect 507397 434088 507469 434144
rect 507397 434054 507416 434088
rect 507450 434054 507469 434088
rect 507397 433998 507469 434054
rect 507397 433964 507416 433998
rect 507450 433964 507469 433998
rect 507397 433908 507469 433964
rect 507397 433874 507416 433908
rect 507450 433874 507469 433908
rect 507397 433818 507469 433874
rect 507397 433784 507416 433818
rect 507450 433784 507469 433818
rect 507397 433728 507469 433784
rect 507397 433694 507416 433728
rect 507450 433694 507469 433728
rect 507397 433638 507469 433694
rect 507397 433604 507416 433638
rect 507450 433604 507469 433638
rect 508287 434290 508306 434324
rect 508340 434290 508359 434324
rect 508287 434234 508359 434290
rect 508287 434200 508306 434234
rect 508340 434200 508359 434234
rect 508287 434144 508359 434200
rect 508287 434110 508306 434144
rect 508340 434110 508359 434144
rect 508287 434054 508359 434110
rect 508287 434020 508306 434054
rect 508340 434020 508359 434054
rect 508287 433964 508359 434020
rect 508287 433930 508306 433964
rect 508340 433930 508359 433964
rect 508287 433874 508359 433930
rect 508287 433840 508306 433874
rect 508340 433840 508359 433874
rect 508287 433784 508359 433840
rect 508287 433750 508306 433784
rect 508340 433750 508359 433784
rect 508287 433694 508359 433750
rect 508287 433660 508306 433694
rect 508340 433660 508359 433694
rect 507397 433565 507469 433604
rect 508287 433604 508359 433660
rect 508287 433570 508306 433604
rect 508340 433570 508359 433604
rect 508287 433565 508359 433570
rect 507397 433546 508359 433565
rect 507397 433512 507510 433546
rect 507544 433512 507600 433546
rect 507634 433512 507690 433546
rect 507724 433512 507780 433546
rect 507814 433512 507870 433546
rect 507904 433512 507960 433546
rect 507994 433512 508050 433546
rect 508084 433512 508140 433546
rect 508174 433512 508230 433546
rect 508264 433512 508359 433546
rect 507397 433493 508359 433512
rect 508685 434436 509647 434455
rect 508685 434402 508817 434436
rect 508851 434402 508907 434436
rect 508941 434402 508997 434436
rect 509031 434402 509087 434436
rect 509121 434402 509177 434436
rect 509211 434402 509267 434436
rect 509301 434402 509357 434436
rect 509391 434402 509447 434436
rect 509481 434402 509537 434436
rect 509571 434402 509647 434436
rect 508685 434383 509647 434402
rect 508685 434358 508757 434383
rect 508685 434324 508704 434358
rect 508738 434324 508757 434358
rect 508685 434268 508757 434324
rect 509575 434324 509647 434383
rect 508685 434234 508704 434268
rect 508738 434234 508757 434268
rect 508685 434178 508757 434234
rect 508685 434144 508704 434178
rect 508738 434144 508757 434178
rect 508685 434088 508757 434144
rect 508685 434054 508704 434088
rect 508738 434054 508757 434088
rect 508685 433998 508757 434054
rect 508685 433964 508704 433998
rect 508738 433964 508757 433998
rect 508685 433908 508757 433964
rect 508685 433874 508704 433908
rect 508738 433874 508757 433908
rect 508685 433818 508757 433874
rect 508685 433784 508704 433818
rect 508738 433784 508757 433818
rect 508685 433728 508757 433784
rect 508685 433694 508704 433728
rect 508738 433694 508757 433728
rect 508685 433638 508757 433694
rect 508685 433604 508704 433638
rect 508738 433604 508757 433638
rect 509575 434290 509594 434324
rect 509628 434290 509647 434324
rect 509575 434234 509647 434290
rect 509575 434200 509594 434234
rect 509628 434200 509647 434234
rect 509575 434144 509647 434200
rect 509575 434110 509594 434144
rect 509628 434110 509647 434144
rect 509575 434054 509647 434110
rect 509575 434020 509594 434054
rect 509628 434020 509647 434054
rect 509575 433964 509647 434020
rect 509575 433930 509594 433964
rect 509628 433930 509647 433964
rect 509575 433874 509647 433930
rect 509575 433840 509594 433874
rect 509628 433840 509647 433874
rect 509575 433784 509647 433840
rect 509575 433750 509594 433784
rect 509628 433750 509647 433784
rect 509575 433694 509647 433750
rect 509575 433660 509594 433694
rect 509628 433660 509647 433694
rect 508685 433565 508757 433604
rect 509575 433604 509647 433660
rect 509575 433570 509594 433604
rect 509628 433570 509647 433604
rect 509575 433565 509647 433570
rect 508685 433546 509647 433565
rect 508685 433512 508798 433546
rect 508832 433512 508888 433546
rect 508922 433512 508978 433546
rect 509012 433512 509068 433546
rect 509102 433512 509158 433546
rect 509192 433512 509248 433546
rect 509282 433512 509338 433546
rect 509372 433512 509428 433546
rect 509462 433512 509518 433546
rect 509552 433512 509647 433546
rect 508685 433493 509647 433512
rect 509973 434436 510935 434455
rect 509973 434402 510105 434436
rect 510139 434402 510195 434436
rect 510229 434402 510285 434436
rect 510319 434402 510375 434436
rect 510409 434402 510465 434436
rect 510499 434402 510555 434436
rect 510589 434402 510645 434436
rect 510679 434402 510735 434436
rect 510769 434402 510825 434436
rect 510859 434402 510935 434436
rect 509973 434383 510935 434402
rect 509973 434358 510045 434383
rect 509973 434324 509992 434358
rect 510026 434324 510045 434358
rect 509973 434268 510045 434324
rect 510863 434324 510935 434383
rect 509973 434234 509992 434268
rect 510026 434234 510045 434268
rect 509973 434178 510045 434234
rect 509973 434144 509992 434178
rect 510026 434144 510045 434178
rect 509973 434088 510045 434144
rect 509973 434054 509992 434088
rect 510026 434054 510045 434088
rect 509973 433998 510045 434054
rect 509973 433964 509992 433998
rect 510026 433964 510045 433998
rect 509973 433908 510045 433964
rect 509973 433874 509992 433908
rect 510026 433874 510045 433908
rect 509973 433818 510045 433874
rect 509973 433784 509992 433818
rect 510026 433784 510045 433818
rect 509973 433728 510045 433784
rect 509973 433694 509992 433728
rect 510026 433694 510045 433728
rect 509973 433638 510045 433694
rect 509973 433604 509992 433638
rect 510026 433604 510045 433638
rect 510863 434290 510882 434324
rect 510916 434290 510935 434324
rect 510863 434234 510935 434290
rect 510863 434200 510882 434234
rect 510916 434200 510935 434234
rect 510863 434144 510935 434200
rect 510863 434110 510882 434144
rect 510916 434110 510935 434144
rect 510863 434054 510935 434110
rect 510863 434020 510882 434054
rect 510916 434020 510935 434054
rect 510863 433964 510935 434020
rect 510863 433930 510882 433964
rect 510916 433930 510935 433964
rect 510863 433874 510935 433930
rect 510863 433840 510882 433874
rect 510916 433840 510935 433874
rect 510863 433784 510935 433840
rect 510863 433750 510882 433784
rect 510916 433750 510935 433784
rect 510863 433694 510935 433750
rect 510863 433660 510882 433694
rect 510916 433660 510935 433694
rect 509973 433565 510045 433604
rect 510863 433604 510935 433660
rect 510863 433570 510882 433604
rect 510916 433570 510935 433604
rect 510863 433565 510935 433570
rect 509973 433546 510935 433565
rect 509973 433512 510086 433546
rect 510120 433512 510176 433546
rect 510210 433512 510266 433546
rect 510300 433512 510356 433546
rect 510390 433512 510446 433546
rect 510480 433512 510536 433546
rect 510570 433512 510626 433546
rect 510660 433512 510716 433546
rect 510750 433512 510806 433546
rect 510840 433512 510935 433546
rect 509973 433493 510935 433512
rect 511261 434436 512223 434455
rect 511261 434402 511393 434436
rect 511427 434402 511483 434436
rect 511517 434402 511573 434436
rect 511607 434402 511663 434436
rect 511697 434402 511753 434436
rect 511787 434402 511843 434436
rect 511877 434402 511933 434436
rect 511967 434402 512023 434436
rect 512057 434402 512113 434436
rect 512147 434402 512223 434436
rect 511261 434383 512223 434402
rect 511261 434358 511333 434383
rect 511261 434324 511280 434358
rect 511314 434324 511333 434358
rect 511261 434268 511333 434324
rect 512151 434324 512223 434383
rect 511261 434234 511280 434268
rect 511314 434234 511333 434268
rect 511261 434178 511333 434234
rect 511261 434144 511280 434178
rect 511314 434144 511333 434178
rect 511261 434088 511333 434144
rect 511261 434054 511280 434088
rect 511314 434054 511333 434088
rect 511261 433998 511333 434054
rect 511261 433964 511280 433998
rect 511314 433964 511333 433998
rect 511261 433908 511333 433964
rect 511261 433874 511280 433908
rect 511314 433874 511333 433908
rect 511261 433818 511333 433874
rect 511261 433784 511280 433818
rect 511314 433784 511333 433818
rect 511261 433728 511333 433784
rect 511261 433694 511280 433728
rect 511314 433694 511333 433728
rect 511261 433638 511333 433694
rect 511261 433604 511280 433638
rect 511314 433604 511333 433638
rect 512151 434290 512170 434324
rect 512204 434290 512223 434324
rect 512151 434234 512223 434290
rect 512151 434200 512170 434234
rect 512204 434200 512223 434234
rect 512151 434144 512223 434200
rect 512151 434110 512170 434144
rect 512204 434110 512223 434144
rect 512151 434054 512223 434110
rect 512151 434020 512170 434054
rect 512204 434020 512223 434054
rect 512151 433964 512223 434020
rect 512151 433930 512170 433964
rect 512204 433930 512223 433964
rect 512151 433874 512223 433930
rect 512151 433840 512170 433874
rect 512204 433840 512223 433874
rect 512151 433784 512223 433840
rect 512151 433750 512170 433784
rect 512204 433750 512223 433784
rect 512151 433694 512223 433750
rect 512151 433660 512170 433694
rect 512204 433660 512223 433694
rect 511261 433565 511333 433604
rect 512151 433604 512223 433660
rect 512151 433570 512170 433604
rect 512204 433570 512223 433604
rect 512151 433565 512223 433570
rect 511261 433546 512223 433565
rect 511261 433512 511374 433546
rect 511408 433512 511464 433546
rect 511498 433512 511554 433546
rect 511588 433512 511644 433546
rect 511678 433512 511734 433546
rect 511768 433512 511824 433546
rect 511858 433512 511914 433546
rect 511948 433512 512004 433546
rect 512038 433512 512094 433546
rect 512128 433512 512223 433546
rect 511261 433493 512223 433512
rect 512549 434436 513511 434455
rect 512549 434402 512681 434436
rect 512715 434402 512771 434436
rect 512805 434402 512861 434436
rect 512895 434402 512951 434436
rect 512985 434402 513041 434436
rect 513075 434402 513131 434436
rect 513165 434402 513221 434436
rect 513255 434402 513311 434436
rect 513345 434402 513401 434436
rect 513435 434402 513511 434436
rect 512549 434383 513511 434402
rect 512549 434358 512621 434383
rect 512549 434324 512568 434358
rect 512602 434324 512621 434358
rect 512549 434268 512621 434324
rect 513439 434324 513511 434383
rect 512549 434234 512568 434268
rect 512602 434234 512621 434268
rect 512549 434178 512621 434234
rect 512549 434144 512568 434178
rect 512602 434144 512621 434178
rect 512549 434088 512621 434144
rect 512549 434054 512568 434088
rect 512602 434054 512621 434088
rect 512549 433998 512621 434054
rect 512549 433964 512568 433998
rect 512602 433964 512621 433998
rect 512549 433908 512621 433964
rect 512549 433874 512568 433908
rect 512602 433874 512621 433908
rect 512549 433818 512621 433874
rect 512549 433784 512568 433818
rect 512602 433784 512621 433818
rect 512549 433728 512621 433784
rect 512549 433694 512568 433728
rect 512602 433694 512621 433728
rect 512549 433638 512621 433694
rect 512549 433604 512568 433638
rect 512602 433604 512621 433638
rect 513439 434290 513458 434324
rect 513492 434290 513511 434324
rect 513439 434234 513511 434290
rect 513439 434200 513458 434234
rect 513492 434200 513511 434234
rect 513439 434144 513511 434200
rect 513439 434110 513458 434144
rect 513492 434110 513511 434144
rect 513439 434054 513511 434110
rect 513439 434020 513458 434054
rect 513492 434020 513511 434054
rect 513439 433964 513511 434020
rect 513439 433930 513458 433964
rect 513492 433930 513511 433964
rect 513439 433874 513511 433930
rect 513439 433840 513458 433874
rect 513492 433840 513511 433874
rect 513439 433784 513511 433840
rect 513439 433750 513458 433784
rect 513492 433750 513511 433784
rect 513439 433694 513511 433750
rect 513439 433660 513458 433694
rect 513492 433660 513511 433694
rect 512549 433565 512621 433604
rect 513439 433604 513511 433660
rect 513439 433570 513458 433604
rect 513492 433570 513511 433604
rect 513439 433565 513511 433570
rect 512549 433546 513511 433565
rect 512549 433512 512662 433546
rect 512696 433512 512752 433546
rect 512786 433512 512842 433546
rect 512876 433512 512932 433546
rect 512966 433512 513022 433546
rect 513056 433512 513112 433546
rect 513146 433512 513202 433546
rect 513236 433512 513292 433546
rect 513326 433512 513382 433546
rect 513416 433512 513511 433546
rect 512549 433493 513511 433512
rect 503533 433148 504495 433167
rect 503533 433114 503665 433148
rect 503699 433114 503755 433148
rect 503789 433114 503845 433148
rect 503879 433114 503935 433148
rect 503969 433114 504025 433148
rect 504059 433114 504115 433148
rect 504149 433114 504205 433148
rect 504239 433114 504295 433148
rect 504329 433114 504385 433148
rect 504419 433114 504495 433148
rect 503533 433095 504495 433114
rect 503533 433070 503605 433095
rect 503533 433036 503552 433070
rect 503586 433036 503605 433070
rect 503533 432980 503605 433036
rect 504423 433036 504495 433095
rect 503533 432946 503552 432980
rect 503586 432946 503605 432980
rect 503533 432890 503605 432946
rect 503533 432856 503552 432890
rect 503586 432856 503605 432890
rect 503533 432800 503605 432856
rect 503533 432766 503552 432800
rect 503586 432766 503605 432800
rect 503533 432710 503605 432766
rect 503533 432676 503552 432710
rect 503586 432676 503605 432710
rect 503533 432620 503605 432676
rect 503533 432586 503552 432620
rect 503586 432586 503605 432620
rect 503533 432530 503605 432586
rect 503533 432496 503552 432530
rect 503586 432496 503605 432530
rect 503533 432440 503605 432496
rect 503533 432406 503552 432440
rect 503586 432406 503605 432440
rect 503533 432350 503605 432406
rect 503533 432316 503552 432350
rect 503586 432316 503605 432350
rect 504423 433002 504442 433036
rect 504476 433002 504495 433036
rect 504423 432946 504495 433002
rect 504423 432912 504442 432946
rect 504476 432912 504495 432946
rect 504423 432856 504495 432912
rect 504423 432822 504442 432856
rect 504476 432822 504495 432856
rect 504423 432766 504495 432822
rect 504423 432732 504442 432766
rect 504476 432732 504495 432766
rect 504423 432676 504495 432732
rect 504423 432642 504442 432676
rect 504476 432642 504495 432676
rect 504423 432586 504495 432642
rect 504423 432552 504442 432586
rect 504476 432552 504495 432586
rect 504423 432496 504495 432552
rect 504423 432462 504442 432496
rect 504476 432462 504495 432496
rect 504423 432406 504495 432462
rect 504423 432372 504442 432406
rect 504476 432372 504495 432406
rect 503533 432277 503605 432316
rect 504423 432316 504495 432372
rect 504423 432282 504442 432316
rect 504476 432282 504495 432316
rect 504423 432277 504495 432282
rect 503533 432258 504495 432277
rect 503533 432224 503646 432258
rect 503680 432224 503736 432258
rect 503770 432224 503826 432258
rect 503860 432224 503916 432258
rect 503950 432224 504006 432258
rect 504040 432224 504096 432258
rect 504130 432224 504186 432258
rect 504220 432224 504276 432258
rect 504310 432224 504366 432258
rect 504400 432224 504495 432258
rect 503533 432205 504495 432224
rect 504821 433148 505783 433167
rect 504821 433114 504953 433148
rect 504987 433114 505043 433148
rect 505077 433114 505133 433148
rect 505167 433114 505223 433148
rect 505257 433114 505313 433148
rect 505347 433114 505403 433148
rect 505437 433114 505493 433148
rect 505527 433114 505583 433148
rect 505617 433114 505673 433148
rect 505707 433114 505783 433148
rect 504821 433095 505783 433114
rect 504821 433070 504893 433095
rect 504821 433036 504840 433070
rect 504874 433036 504893 433070
rect 504821 432980 504893 433036
rect 505711 433036 505783 433095
rect 504821 432946 504840 432980
rect 504874 432946 504893 432980
rect 504821 432890 504893 432946
rect 504821 432856 504840 432890
rect 504874 432856 504893 432890
rect 504821 432800 504893 432856
rect 504821 432766 504840 432800
rect 504874 432766 504893 432800
rect 504821 432710 504893 432766
rect 504821 432676 504840 432710
rect 504874 432676 504893 432710
rect 504821 432620 504893 432676
rect 504821 432586 504840 432620
rect 504874 432586 504893 432620
rect 504821 432530 504893 432586
rect 504821 432496 504840 432530
rect 504874 432496 504893 432530
rect 504821 432440 504893 432496
rect 504821 432406 504840 432440
rect 504874 432406 504893 432440
rect 504821 432350 504893 432406
rect 504821 432316 504840 432350
rect 504874 432316 504893 432350
rect 505711 433002 505730 433036
rect 505764 433002 505783 433036
rect 505711 432946 505783 433002
rect 505711 432912 505730 432946
rect 505764 432912 505783 432946
rect 505711 432856 505783 432912
rect 505711 432822 505730 432856
rect 505764 432822 505783 432856
rect 505711 432766 505783 432822
rect 505711 432732 505730 432766
rect 505764 432732 505783 432766
rect 505711 432676 505783 432732
rect 505711 432642 505730 432676
rect 505764 432642 505783 432676
rect 505711 432586 505783 432642
rect 505711 432552 505730 432586
rect 505764 432552 505783 432586
rect 505711 432496 505783 432552
rect 505711 432462 505730 432496
rect 505764 432462 505783 432496
rect 505711 432406 505783 432462
rect 505711 432372 505730 432406
rect 505764 432372 505783 432406
rect 504821 432277 504893 432316
rect 505711 432316 505783 432372
rect 505711 432282 505730 432316
rect 505764 432282 505783 432316
rect 505711 432277 505783 432282
rect 504821 432258 505783 432277
rect 504821 432224 504934 432258
rect 504968 432224 505024 432258
rect 505058 432224 505114 432258
rect 505148 432224 505204 432258
rect 505238 432224 505294 432258
rect 505328 432224 505384 432258
rect 505418 432224 505474 432258
rect 505508 432224 505564 432258
rect 505598 432224 505654 432258
rect 505688 432224 505783 432258
rect 504821 432205 505783 432224
rect 506109 433148 507071 433167
rect 506109 433114 506241 433148
rect 506275 433114 506331 433148
rect 506365 433114 506421 433148
rect 506455 433114 506511 433148
rect 506545 433114 506601 433148
rect 506635 433114 506691 433148
rect 506725 433114 506781 433148
rect 506815 433114 506871 433148
rect 506905 433114 506961 433148
rect 506995 433114 507071 433148
rect 506109 433095 507071 433114
rect 506109 433070 506181 433095
rect 506109 433036 506128 433070
rect 506162 433036 506181 433070
rect 506109 432980 506181 433036
rect 506999 433036 507071 433095
rect 506109 432946 506128 432980
rect 506162 432946 506181 432980
rect 506109 432890 506181 432946
rect 506109 432856 506128 432890
rect 506162 432856 506181 432890
rect 506109 432800 506181 432856
rect 506109 432766 506128 432800
rect 506162 432766 506181 432800
rect 506109 432710 506181 432766
rect 506109 432676 506128 432710
rect 506162 432676 506181 432710
rect 506109 432620 506181 432676
rect 506109 432586 506128 432620
rect 506162 432586 506181 432620
rect 506109 432530 506181 432586
rect 506109 432496 506128 432530
rect 506162 432496 506181 432530
rect 506109 432440 506181 432496
rect 506109 432406 506128 432440
rect 506162 432406 506181 432440
rect 506109 432350 506181 432406
rect 506109 432316 506128 432350
rect 506162 432316 506181 432350
rect 506999 433002 507018 433036
rect 507052 433002 507071 433036
rect 506999 432946 507071 433002
rect 506999 432912 507018 432946
rect 507052 432912 507071 432946
rect 506999 432856 507071 432912
rect 506999 432822 507018 432856
rect 507052 432822 507071 432856
rect 506999 432766 507071 432822
rect 506999 432732 507018 432766
rect 507052 432732 507071 432766
rect 506999 432676 507071 432732
rect 506999 432642 507018 432676
rect 507052 432642 507071 432676
rect 506999 432586 507071 432642
rect 506999 432552 507018 432586
rect 507052 432552 507071 432586
rect 506999 432496 507071 432552
rect 506999 432462 507018 432496
rect 507052 432462 507071 432496
rect 506999 432406 507071 432462
rect 506999 432372 507018 432406
rect 507052 432372 507071 432406
rect 506109 432277 506181 432316
rect 506999 432316 507071 432372
rect 506999 432282 507018 432316
rect 507052 432282 507071 432316
rect 506999 432277 507071 432282
rect 506109 432258 507071 432277
rect 506109 432224 506222 432258
rect 506256 432224 506312 432258
rect 506346 432224 506402 432258
rect 506436 432224 506492 432258
rect 506526 432224 506582 432258
rect 506616 432224 506672 432258
rect 506706 432224 506762 432258
rect 506796 432224 506852 432258
rect 506886 432224 506942 432258
rect 506976 432224 507071 432258
rect 506109 432205 507071 432224
rect 507397 433148 508359 433167
rect 507397 433114 507529 433148
rect 507563 433114 507619 433148
rect 507653 433114 507709 433148
rect 507743 433114 507799 433148
rect 507833 433114 507889 433148
rect 507923 433114 507979 433148
rect 508013 433114 508069 433148
rect 508103 433114 508159 433148
rect 508193 433114 508249 433148
rect 508283 433114 508359 433148
rect 507397 433095 508359 433114
rect 507397 433070 507469 433095
rect 507397 433036 507416 433070
rect 507450 433036 507469 433070
rect 507397 432980 507469 433036
rect 508287 433036 508359 433095
rect 507397 432946 507416 432980
rect 507450 432946 507469 432980
rect 507397 432890 507469 432946
rect 507397 432856 507416 432890
rect 507450 432856 507469 432890
rect 507397 432800 507469 432856
rect 507397 432766 507416 432800
rect 507450 432766 507469 432800
rect 507397 432710 507469 432766
rect 507397 432676 507416 432710
rect 507450 432676 507469 432710
rect 507397 432620 507469 432676
rect 507397 432586 507416 432620
rect 507450 432586 507469 432620
rect 507397 432530 507469 432586
rect 507397 432496 507416 432530
rect 507450 432496 507469 432530
rect 507397 432440 507469 432496
rect 507397 432406 507416 432440
rect 507450 432406 507469 432440
rect 507397 432350 507469 432406
rect 507397 432316 507416 432350
rect 507450 432316 507469 432350
rect 508287 433002 508306 433036
rect 508340 433002 508359 433036
rect 508287 432946 508359 433002
rect 508287 432912 508306 432946
rect 508340 432912 508359 432946
rect 508287 432856 508359 432912
rect 508287 432822 508306 432856
rect 508340 432822 508359 432856
rect 508287 432766 508359 432822
rect 508287 432732 508306 432766
rect 508340 432732 508359 432766
rect 508287 432676 508359 432732
rect 508287 432642 508306 432676
rect 508340 432642 508359 432676
rect 508287 432586 508359 432642
rect 508287 432552 508306 432586
rect 508340 432552 508359 432586
rect 508287 432496 508359 432552
rect 508287 432462 508306 432496
rect 508340 432462 508359 432496
rect 508287 432406 508359 432462
rect 508287 432372 508306 432406
rect 508340 432372 508359 432406
rect 507397 432277 507469 432316
rect 508287 432316 508359 432372
rect 508287 432282 508306 432316
rect 508340 432282 508359 432316
rect 508287 432277 508359 432282
rect 507397 432258 508359 432277
rect 507397 432224 507510 432258
rect 507544 432224 507600 432258
rect 507634 432224 507690 432258
rect 507724 432224 507780 432258
rect 507814 432224 507870 432258
rect 507904 432224 507960 432258
rect 507994 432224 508050 432258
rect 508084 432224 508140 432258
rect 508174 432224 508230 432258
rect 508264 432224 508359 432258
rect 507397 432205 508359 432224
rect 508685 433148 509647 433167
rect 508685 433114 508817 433148
rect 508851 433114 508907 433148
rect 508941 433114 508997 433148
rect 509031 433114 509087 433148
rect 509121 433114 509177 433148
rect 509211 433114 509267 433148
rect 509301 433114 509357 433148
rect 509391 433114 509447 433148
rect 509481 433114 509537 433148
rect 509571 433114 509647 433148
rect 508685 433095 509647 433114
rect 508685 433070 508757 433095
rect 508685 433036 508704 433070
rect 508738 433036 508757 433070
rect 508685 432980 508757 433036
rect 509575 433036 509647 433095
rect 508685 432946 508704 432980
rect 508738 432946 508757 432980
rect 508685 432890 508757 432946
rect 508685 432856 508704 432890
rect 508738 432856 508757 432890
rect 508685 432800 508757 432856
rect 508685 432766 508704 432800
rect 508738 432766 508757 432800
rect 508685 432710 508757 432766
rect 508685 432676 508704 432710
rect 508738 432676 508757 432710
rect 508685 432620 508757 432676
rect 508685 432586 508704 432620
rect 508738 432586 508757 432620
rect 508685 432530 508757 432586
rect 508685 432496 508704 432530
rect 508738 432496 508757 432530
rect 508685 432440 508757 432496
rect 508685 432406 508704 432440
rect 508738 432406 508757 432440
rect 508685 432350 508757 432406
rect 508685 432316 508704 432350
rect 508738 432316 508757 432350
rect 509575 433002 509594 433036
rect 509628 433002 509647 433036
rect 509575 432946 509647 433002
rect 509575 432912 509594 432946
rect 509628 432912 509647 432946
rect 509575 432856 509647 432912
rect 509575 432822 509594 432856
rect 509628 432822 509647 432856
rect 509575 432766 509647 432822
rect 509575 432732 509594 432766
rect 509628 432732 509647 432766
rect 509575 432676 509647 432732
rect 509575 432642 509594 432676
rect 509628 432642 509647 432676
rect 509575 432586 509647 432642
rect 509575 432552 509594 432586
rect 509628 432552 509647 432586
rect 509575 432496 509647 432552
rect 509575 432462 509594 432496
rect 509628 432462 509647 432496
rect 509575 432406 509647 432462
rect 509575 432372 509594 432406
rect 509628 432372 509647 432406
rect 508685 432277 508757 432316
rect 509575 432316 509647 432372
rect 509575 432282 509594 432316
rect 509628 432282 509647 432316
rect 509575 432277 509647 432282
rect 508685 432258 509647 432277
rect 508685 432224 508798 432258
rect 508832 432224 508888 432258
rect 508922 432224 508978 432258
rect 509012 432224 509068 432258
rect 509102 432224 509158 432258
rect 509192 432224 509248 432258
rect 509282 432224 509338 432258
rect 509372 432224 509428 432258
rect 509462 432224 509518 432258
rect 509552 432224 509647 432258
rect 508685 432205 509647 432224
rect 509973 433148 510935 433167
rect 509973 433114 510105 433148
rect 510139 433114 510195 433148
rect 510229 433114 510285 433148
rect 510319 433114 510375 433148
rect 510409 433114 510465 433148
rect 510499 433114 510555 433148
rect 510589 433114 510645 433148
rect 510679 433114 510735 433148
rect 510769 433114 510825 433148
rect 510859 433114 510935 433148
rect 509973 433095 510935 433114
rect 509973 433070 510045 433095
rect 509973 433036 509992 433070
rect 510026 433036 510045 433070
rect 509973 432980 510045 433036
rect 510863 433036 510935 433095
rect 509973 432946 509992 432980
rect 510026 432946 510045 432980
rect 509973 432890 510045 432946
rect 509973 432856 509992 432890
rect 510026 432856 510045 432890
rect 509973 432800 510045 432856
rect 509973 432766 509992 432800
rect 510026 432766 510045 432800
rect 509973 432710 510045 432766
rect 509973 432676 509992 432710
rect 510026 432676 510045 432710
rect 509973 432620 510045 432676
rect 509973 432586 509992 432620
rect 510026 432586 510045 432620
rect 509973 432530 510045 432586
rect 509973 432496 509992 432530
rect 510026 432496 510045 432530
rect 509973 432440 510045 432496
rect 509973 432406 509992 432440
rect 510026 432406 510045 432440
rect 509973 432350 510045 432406
rect 509973 432316 509992 432350
rect 510026 432316 510045 432350
rect 510863 433002 510882 433036
rect 510916 433002 510935 433036
rect 510863 432946 510935 433002
rect 510863 432912 510882 432946
rect 510916 432912 510935 432946
rect 510863 432856 510935 432912
rect 510863 432822 510882 432856
rect 510916 432822 510935 432856
rect 510863 432766 510935 432822
rect 510863 432732 510882 432766
rect 510916 432732 510935 432766
rect 510863 432676 510935 432732
rect 510863 432642 510882 432676
rect 510916 432642 510935 432676
rect 510863 432586 510935 432642
rect 510863 432552 510882 432586
rect 510916 432552 510935 432586
rect 510863 432496 510935 432552
rect 510863 432462 510882 432496
rect 510916 432462 510935 432496
rect 510863 432406 510935 432462
rect 510863 432372 510882 432406
rect 510916 432372 510935 432406
rect 509973 432277 510045 432316
rect 510863 432316 510935 432372
rect 510863 432282 510882 432316
rect 510916 432282 510935 432316
rect 510863 432277 510935 432282
rect 509973 432258 510935 432277
rect 509973 432224 510086 432258
rect 510120 432224 510176 432258
rect 510210 432224 510266 432258
rect 510300 432224 510356 432258
rect 510390 432224 510446 432258
rect 510480 432224 510536 432258
rect 510570 432224 510626 432258
rect 510660 432224 510716 432258
rect 510750 432224 510806 432258
rect 510840 432224 510935 432258
rect 509973 432205 510935 432224
rect 511261 433148 512223 433167
rect 511261 433114 511393 433148
rect 511427 433114 511483 433148
rect 511517 433114 511573 433148
rect 511607 433114 511663 433148
rect 511697 433114 511753 433148
rect 511787 433114 511843 433148
rect 511877 433114 511933 433148
rect 511967 433114 512023 433148
rect 512057 433114 512113 433148
rect 512147 433114 512223 433148
rect 511261 433095 512223 433114
rect 511261 433070 511333 433095
rect 511261 433036 511280 433070
rect 511314 433036 511333 433070
rect 511261 432980 511333 433036
rect 512151 433036 512223 433095
rect 511261 432946 511280 432980
rect 511314 432946 511333 432980
rect 511261 432890 511333 432946
rect 511261 432856 511280 432890
rect 511314 432856 511333 432890
rect 511261 432800 511333 432856
rect 511261 432766 511280 432800
rect 511314 432766 511333 432800
rect 511261 432710 511333 432766
rect 511261 432676 511280 432710
rect 511314 432676 511333 432710
rect 511261 432620 511333 432676
rect 511261 432586 511280 432620
rect 511314 432586 511333 432620
rect 511261 432530 511333 432586
rect 511261 432496 511280 432530
rect 511314 432496 511333 432530
rect 511261 432440 511333 432496
rect 511261 432406 511280 432440
rect 511314 432406 511333 432440
rect 511261 432350 511333 432406
rect 511261 432316 511280 432350
rect 511314 432316 511333 432350
rect 512151 433002 512170 433036
rect 512204 433002 512223 433036
rect 512151 432946 512223 433002
rect 512151 432912 512170 432946
rect 512204 432912 512223 432946
rect 512151 432856 512223 432912
rect 512151 432822 512170 432856
rect 512204 432822 512223 432856
rect 512151 432766 512223 432822
rect 512151 432732 512170 432766
rect 512204 432732 512223 432766
rect 512151 432676 512223 432732
rect 512151 432642 512170 432676
rect 512204 432642 512223 432676
rect 512151 432586 512223 432642
rect 512151 432552 512170 432586
rect 512204 432552 512223 432586
rect 512151 432496 512223 432552
rect 512151 432462 512170 432496
rect 512204 432462 512223 432496
rect 512151 432406 512223 432462
rect 512151 432372 512170 432406
rect 512204 432372 512223 432406
rect 511261 432277 511333 432316
rect 512151 432316 512223 432372
rect 512151 432282 512170 432316
rect 512204 432282 512223 432316
rect 512151 432277 512223 432282
rect 511261 432258 512223 432277
rect 511261 432224 511374 432258
rect 511408 432224 511464 432258
rect 511498 432224 511554 432258
rect 511588 432224 511644 432258
rect 511678 432224 511734 432258
rect 511768 432224 511824 432258
rect 511858 432224 511914 432258
rect 511948 432224 512004 432258
rect 512038 432224 512094 432258
rect 512128 432224 512223 432258
rect 511261 432205 512223 432224
rect 512549 433148 513511 433167
rect 512549 433114 512681 433148
rect 512715 433114 512771 433148
rect 512805 433114 512861 433148
rect 512895 433114 512951 433148
rect 512985 433114 513041 433148
rect 513075 433114 513131 433148
rect 513165 433114 513221 433148
rect 513255 433114 513311 433148
rect 513345 433114 513401 433148
rect 513435 433114 513511 433148
rect 512549 433095 513511 433114
rect 512549 433070 512621 433095
rect 512549 433036 512568 433070
rect 512602 433036 512621 433070
rect 512549 432980 512621 433036
rect 513439 433036 513511 433095
rect 512549 432946 512568 432980
rect 512602 432946 512621 432980
rect 512549 432890 512621 432946
rect 512549 432856 512568 432890
rect 512602 432856 512621 432890
rect 512549 432800 512621 432856
rect 512549 432766 512568 432800
rect 512602 432766 512621 432800
rect 512549 432710 512621 432766
rect 512549 432676 512568 432710
rect 512602 432676 512621 432710
rect 512549 432620 512621 432676
rect 512549 432586 512568 432620
rect 512602 432586 512621 432620
rect 512549 432530 512621 432586
rect 512549 432496 512568 432530
rect 512602 432496 512621 432530
rect 512549 432440 512621 432496
rect 512549 432406 512568 432440
rect 512602 432406 512621 432440
rect 512549 432350 512621 432406
rect 512549 432316 512568 432350
rect 512602 432316 512621 432350
rect 513439 433002 513458 433036
rect 513492 433002 513511 433036
rect 513439 432946 513511 433002
rect 513439 432912 513458 432946
rect 513492 432912 513511 432946
rect 513439 432856 513511 432912
rect 513439 432822 513458 432856
rect 513492 432822 513511 432856
rect 513439 432766 513511 432822
rect 513439 432732 513458 432766
rect 513492 432732 513511 432766
rect 513439 432676 513511 432732
rect 513439 432642 513458 432676
rect 513492 432642 513511 432676
rect 513439 432586 513511 432642
rect 513439 432552 513458 432586
rect 513492 432552 513511 432586
rect 513439 432496 513511 432552
rect 513439 432462 513458 432496
rect 513492 432462 513511 432496
rect 513439 432406 513511 432462
rect 513439 432372 513458 432406
rect 513492 432372 513511 432406
rect 512549 432277 512621 432316
rect 513439 432316 513511 432372
rect 513439 432282 513458 432316
rect 513492 432282 513511 432316
rect 513439 432277 513511 432282
rect 512549 432258 513511 432277
rect 512549 432224 512662 432258
rect 512696 432224 512752 432258
rect 512786 432224 512842 432258
rect 512876 432224 512932 432258
rect 512966 432224 513022 432258
rect 513056 432224 513112 432258
rect 513146 432224 513202 432258
rect 513236 432224 513292 432258
rect 513326 432224 513382 432258
rect 513416 432224 513511 432258
rect 512549 432205 513511 432224
rect 562156 455178 562252 455212
rect 567482 455178 567578 455212
rect 562156 455115 562190 455178
rect 567544 455115 567578 455178
rect 562156 453950 562190 454013
rect 567544 453950 567578 454013
rect 562156 453916 562252 453950
rect 567482 453916 567578 453950
<< psubdiffcont >>
rect 572412 495514 577642 495548
rect 572316 494358 572350 495452
rect 577704 494358 577738 495452
rect 572412 494262 577642 494296
rect 500368 432068 501368 475308
rect 502392 474284 526544 475284
rect 506532 472856 507108 473256
rect 507186 470878 507262 471870
rect 506532 469490 507108 469890
rect 506468 468286 508068 468386
rect 506468 462786 508068 462886
rect 510476 462382 510808 468834
rect 525696 461284 526462 472468
rect 516622 460138 522926 460708
rect 516622 456894 522926 457464
rect 516622 451934 522926 452504
rect 503486 438414 503520 438448
rect 503576 438414 503610 438448
rect 503666 438414 503700 438448
rect 503756 438414 503790 438448
rect 503846 438414 503880 438448
rect 503936 438414 503970 438448
rect 504026 438414 504060 438448
rect 504116 438414 504150 438448
rect 504206 438414 504240 438448
rect 504296 438414 504330 438448
rect 504386 438414 504420 438448
rect 504476 438414 504510 438448
rect 504566 438414 504600 438448
rect 504774 438414 504808 438448
rect 504864 438414 504898 438448
rect 504954 438414 504988 438448
rect 505044 438414 505078 438448
rect 505134 438414 505168 438448
rect 505224 438414 505258 438448
rect 505314 438414 505348 438448
rect 505404 438414 505438 438448
rect 505494 438414 505528 438448
rect 505584 438414 505618 438448
rect 505674 438414 505708 438448
rect 505764 438414 505798 438448
rect 505854 438414 505888 438448
rect 506062 438414 506096 438448
rect 506152 438414 506186 438448
rect 506242 438414 506276 438448
rect 506332 438414 506366 438448
rect 506422 438414 506456 438448
rect 506512 438414 506546 438448
rect 506602 438414 506636 438448
rect 506692 438414 506726 438448
rect 506782 438414 506816 438448
rect 506872 438414 506906 438448
rect 506962 438414 506996 438448
rect 507052 438414 507086 438448
rect 507142 438414 507176 438448
rect 507350 438414 507384 438448
rect 507440 438414 507474 438448
rect 507530 438414 507564 438448
rect 507620 438414 507654 438448
rect 507710 438414 507744 438448
rect 507800 438414 507834 438448
rect 507890 438414 507924 438448
rect 507980 438414 508014 438448
rect 508070 438414 508104 438448
rect 508160 438414 508194 438448
rect 508250 438414 508284 438448
rect 508340 438414 508374 438448
rect 508430 438414 508464 438448
rect 508638 438414 508672 438448
rect 508728 438414 508762 438448
rect 508818 438414 508852 438448
rect 508908 438414 508942 438448
rect 508998 438414 509032 438448
rect 509088 438414 509122 438448
rect 509178 438414 509212 438448
rect 509268 438414 509302 438448
rect 509358 438414 509392 438448
rect 509448 438414 509482 438448
rect 509538 438414 509572 438448
rect 509628 438414 509662 438448
rect 509718 438414 509752 438448
rect 509926 438414 509960 438448
rect 510016 438414 510050 438448
rect 510106 438414 510140 438448
rect 510196 438414 510230 438448
rect 510286 438414 510320 438448
rect 510376 438414 510410 438448
rect 510466 438414 510500 438448
rect 510556 438414 510590 438448
rect 510646 438414 510680 438448
rect 510736 438414 510770 438448
rect 510826 438414 510860 438448
rect 510916 438414 510950 438448
rect 511006 438414 511040 438448
rect 511214 438414 511248 438448
rect 511304 438414 511338 438448
rect 511394 438414 511428 438448
rect 511484 438414 511518 438448
rect 511574 438414 511608 438448
rect 511664 438414 511698 438448
rect 511754 438414 511788 438448
rect 511844 438414 511878 438448
rect 511934 438414 511968 438448
rect 512024 438414 512058 438448
rect 512114 438414 512148 438448
rect 512204 438414 512238 438448
rect 512294 438414 512328 438448
rect 512502 438414 512536 438448
rect 512592 438414 512626 438448
rect 512682 438414 512716 438448
rect 512772 438414 512806 438448
rect 512862 438414 512896 438448
rect 512952 438414 512986 438448
rect 513042 438414 513076 438448
rect 513132 438414 513166 438448
rect 513222 438414 513256 438448
rect 513312 438414 513346 438448
rect 513402 438414 513436 438448
rect 513492 438414 513526 438448
rect 513582 438414 513616 438448
rect 503402 438318 503436 438352
rect 503402 438228 503436 438262
rect 503402 438138 503436 438172
rect 503402 438048 503436 438082
rect 503402 437958 503436 437992
rect 503402 437868 503436 437902
rect 503402 437778 503436 437812
rect 503402 437688 503436 437722
rect 503402 437598 503436 437632
rect 503402 437508 503436 437542
rect 503402 437418 503436 437452
rect 503402 437328 503436 437362
rect 504589 438318 504623 438352
rect 504690 438318 504724 438352
rect 504589 438228 504623 438262
rect 504690 438228 504724 438262
rect 504589 438138 504623 438172
rect 504690 438138 504724 438172
rect 504589 438048 504623 438082
rect 504690 438048 504724 438082
rect 504589 437958 504623 437992
rect 504690 437958 504724 437992
rect 504589 437868 504623 437902
rect 504690 437868 504724 437902
rect 504589 437778 504623 437812
rect 504690 437778 504724 437812
rect 504589 437688 504623 437722
rect 504690 437688 504724 437722
rect 504589 437598 504623 437632
rect 504690 437598 504724 437632
rect 504589 437508 504623 437542
rect 504690 437508 504724 437542
rect 504589 437418 504623 437452
rect 504690 437418 504724 437452
rect 504589 437328 504623 437362
rect 504690 437328 504724 437362
rect 505877 438318 505911 438352
rect 505978 438318 506012 438352
rect 505877 438228 505911 438262
rect 505978 438228 506012 438262
rect 505877 438138 505911 438172
rect 505978 438138 506012 438172
rect 505877 438048 505911 438082
rect 505978 438048 506012 438082
rect 505877 437958 505911 437992
rect 505978 437958 506012 437992
rect 505877 437868 505911 437902
rect 505978 437868 506012 437902
rect 505877 437778 505911 437812
rect 505978 437778 506012 437812
rect 505877 437688 505911 437722
rect 505978 437688 506012 437722
rect 505877 437598 505911 437632
rect 505978 437598 506012 437632
rect 505877 437508 505911 437542
rect 505978 437508 506012 437542
rect 505877 437418 505911 437452
rect 505978 437418 506012 437452
rect 505877 437328 505911 437362
rect 505978 437328 506012 437362
rect 507165 438318 507199 438352
rect 507266 438318 507300 438352
rect 507165 438228 507199 438262
rect 507266 438228 507300 438262
rect 507165 438138 507199 438172
rect 507266 438138 507300 438172
rect 507165 438048 507199 438082
rect 507266 438048 507300 438082
rect 507165 437958 507199 437992
rect 507266 437958 507300 437992
rect 507165 437868 507199 437902
rect 507266 437868 507300 437902
rect 507165 437778 507199 437812
rect 507266 437778 507300 437812
rect 507165 437688 507199 437722
rect 507266 437688 507300 437722
rect 507165 437598 507199 437632
rect 507266 437598 507300 437632
rect 507165 437508 507199 437542
rect 507266 437508 507300 437542
rect 507165 437418 507199 437452
rect 507266 437418 507300 437452
rect 507165 437328 507199 437362
rect 507266 437328 507300 437362
rect 508453 438318 508487 438352
rect 508554 438318 508588 438352
rect 508453 438228 508487 438262
rect 508554 438228 508588 438262
rect 508453 438138 508487 438172
rect 508554 438138 508588 438172
rect 508453 438048 508487 438082
rect 508554 438048 508588 438082
rect 508453 437958 508487 437992
rect 508554 437958 508588 437992
rect 508453 437868 508487 437902
rect 508554 437868 508588 437902
rect 508453 437778 508487 437812
rect 508554 437778 508588 437812
rect 508453 437688 508487 437722
rect 508554 437688 508588 437722
rect 508453 437598 508487 437632
rect 508554 437598 508588 437632
rect 508453 437508 508487 437542
rect 508554 437508 508588 437542
rect 508453 437418 508487 437452
rect 508554 437418 508588 437452
rect 508453 437328 508487 437362
rect 508554 437328 508588 437362
rect 509741 438318 509775 438352
rect 509842 438318 509876 438352
rect 509741 438228 509775 438262
rect 509842 438228 509876 438262
rect 509741 438138 509775 438172
rect 509842 438138 509876 438172
rect 509741 438048 509775 438082
rect 509842 438048 509876 438082
rect 509741 437958 509775 437992
rect 509842 437958 509876 437992
rect 509741 437868 509775 437902
rect 509842 437868 509876 437902
rect 509741 437778 509775 437812
rect 509842 437778 509876 437812
rect 509741 437688 509775 437722
rect 509842 437688 509876 437722
rect 509741 437598 509775 437632
rect 509842 437598 509876 437632
rect 509741 437508 509775 437542
rect 509842 437508 509876 437542
rect 509741 437418 509775 437452
rect 509842 437418 509876 437452
rect 509741 437328 509775 437362
rect 509842 437328 509876 437362
rect 511029 438318 511063 438352
rect 511130 438318 511164 438352
rect 511029 438228 511063 438262
rect 511130 438228 511164 438262
rect 511029 438138 511063 438172
rect 511130 438138 511164 438172
rect 511029 438048 511063 438082
rect 511130 438048 511164 438082
rect 511029 437958 511063 437992
rect 511130 437958 511164 437992
rect 511029 437868 511063 437902
rect 511130 437868 511164 437902
rect 511029 437778 511063 437812
rect 511130 437778 511164 437812
rect 511029 437688 511063 437722
rect 511130 437688 511164 437722
rect 511029 437598 511063 437632
rect 511130 437598 511164 437632
rect 511029 437508 511063 437542
rect 511130 437508 511164 437542
rect 511029 437418 511063 437452
rect 511130 437418 511164 437452
rect 511029 437328 511063 437362
rect 511130 437328 511164 437362
rect 512317 438318 512351 438352
rect 512418 438318 512452 438352
rect 512317 438228 512351 438262
rect 512418 438228 512452 438262
rect 512317 438138 512351 438172
rect 512418 438138 512452 438172
rect 512317 438048 512351 438082
rect 512418 438048 512452 438082
rect 512317 437958 512351 437992
rect 512418 437958 512452 437992
rect 512317 437868 512351 437902
rect 512418 437868 512452 437902
rect 512317 437778 512351 437812
rect 512418 437778 512452 437812
rect 512317 437688 512351 437722
rect 512418 437688 512452 437722
rect 512317 437598 512351 437632
rect 512418 437598 512452 437632
rect 512317 437508 512351 437542
rect 512418 437508 512452 437542
rect 512317 437418 512351 437452
rect 512418 437418 512452 437452
rect 512317 437328 512351 437362
rect 512418 437328 512452 437362
rect 513605 438318 513639 438352
rect 513605 438228 513639 438262
rect 513605 438138 513639 438172
rect 513605 438048 513639 438082
rect 513605 437958 513639 437992
rect 513605 437868 513639 437902
rect 513605 437778 513639 437812
rect 513605 437688 513639 437722
rect 513605 437598 513639 437632
rect 513605 437508 513639 437542
rect 513605 437418 513639 437452
rect 513605 437328 513639 437362
rect 503486 437227 503520 437261
rect 503576 437227 503610 437261
rect 503666 437227 503700 437261
rect 503756 437227 503790 437261
rect 503846 437227 503880 437261
rect 503936 437227 503970 437261
rect 504026 437227 504060 437261
rect 504116 437227 504150 437261
rect 504206 437227 504240 437261
rect 504296 437227 504330 437261
rect 504386 437227 504420 437261
rect 504476 437227 504510 437261
rect 504566 437227 504600 437261
rect 504774 437227 504808 437261
rect 504864 437227 504898 437261
rect 504954 437227 504988 437261
rect 505044 437227 505078 437261
rect 505134 437227 505168 437261
rect 505224 437227 505258 437261
rect 505314 437227 505348 437261
rect 505404 437227 505438 437261
rect 505494 437227 505528 437261
rect 505584 437227 505618 437261
rect 505674 437227 505708 437261
rect 505764 437227 505798 437261
rect 505854 437227 505888 437261
rect 506062 437227 506096 437261
rect 506152 437227 506186 437261
rect 506242 437227 506276 437261
rect 506332 437227 506366 437261
rect 506422 437227 506456 437261
rect 506512 437227 506546 437261
rect 506602 437227 506636 437261
rect 506692 437227 506726 437261
rect 506782 437227 506816 437261
rect 506872 437227 506906 437261
rect 506962 437227 506996 437261
rect 507052 437227 507086 437261
rect 507142 437227 507176 437261
rect 507350 437227 507384 437261
rect 507440 437227 507474 437261
rect 507530 437227 507564 437261
rect 507620 437227 507654 437261
rect 507710 437227 507744 437261
rect 507800 437227 507834 437261
rect 507890 437227 507924 437261
rect 507980 437227 508014 437261
rect 508070 437227 508104 437261
rect 508160 437227 508194 437261
rect 508250 437227 508284 437261
rect 508340 437227 508374 437261
rect 508430 437227 508464 437261
rect 508638 437227 508672 437261
rect 508728 437227 508762 437261
rect 508818 437227 508852 437261
rect 508908 437227 508942 437261
rect 508998 437227 509032 437261
rect 509088 437227 509122 437261
rect 509178 437227 509212 437261
rect 509268 437227 509302 437261
rect 509358 437227 509392 437261
rect 509448 437227 509482 437261
rect 509538 437227 509572 437261
rect 509628 437227 509662 437261
rect 509718 437227 509752 437261
rect 509926 437227 509960 437261
rect 510016 437227 510050 437261
rect 510106 437227 510140 437261
rect 510196 437227 510230 437261
rect 510286 437227 510320 437261
rect 510376 437227 510410 437261
rect 510466 437227 510500 437261
rect 510556 437227 510590 437261
rect 510646 437227 510680 437261
rect 510736 437227 510770 437261
rect 510826 437227 510860 437261
rect 510916 437227 510950 437261
rect 511006 437227 511040 437261
rect 511214 437227 511248 437261
rect 511304 437227 511338 437261
rect 511394 437227 511428 437261
rect 511484 437227 511518 437261
rect 511574 437227 511608 437261
rect 511664 437227 511698 437261
rect 511754 437227 511788 437261
rect 511844 437227 511878 437261
rect 511934 437227 511968 437261
rect 512024 437227 512058 437261
rect 512114 437227 512148 437261
rect 512204 437227 512238 437261
rect 512294 437227 512328 437261
rect 512502 437227 512536 437261
rect 512592 437227 512626 437261
rect 512682 437227 512716 437261
rect 512772 437227 512806 437261
rect 512862 437227 512896 437261
rect 512952 437227 512986 437261
rect 513042 437227 513076 437261
rect 513132 437227 513166 437261
rect 513222 437227 513256 437261
rect 513312 437227 513346 437261
rect 513402 437227 513436 437261
rect 513492 437227 513526 437261
rect 513582 437227 513616 437261
rect 516622 437246 522926 437816
rect 503486 437126 503520 437160
rect 503576 437126 503610 437160
rect 503666 437126 503700 437160
rect 503756 437126 503790 437160
rect 503846 437126 503880 437160
rect 503936 437126 503970 437160
rect 504026 437126 504060 437160
rect 504116 437126 504150 437160
rect 504206 437126 504240 437160
rect 504296 437126 504330 437160
rect 504386 437126 504420 437160
rect 504476 437126 504510 437160
rect 504566 437126 504600 437160
rect 504774 437126 504808 437160
rect 504864 437126 504898 437160
rect 504954 437126 504988 437160
rect 505044 437126 505078 437160
rect 505134 437126 505168 437160
rect 505224 437126 505258 437160
rect 505314 437126 505348 437160
rect 505404 437126 505438 437160
rect 505494 437126 505528 437160
rect 505584 437126 505618 437160
rect 505674 437126 505708 437160
rect 505764 437126 505798 437160
rect 505854 437126 505888 437160
rect 506062 437126 506096 437160
rect 506152 437126 506186 437160
rect 506242 437126 506276 437160
rect 506332 437126 506366 437160
rect 506422 437126 506456 437160
rect 506512 437126 506546 437160
rect 506602 437126 506636 437160
rect 506692 437126 506726 437160
rect 506782 437126 506816 437160
rect 506872 437126 506906 437160
rect 506962 437126 506996 437160
rect 507052 437126 507086 437160
rect 507142 437126 507176 437160
rect 507350 437126 507384 437160
rect 507440 437126 507474 437160
rect 507530 437126 507564 437160
rect 507620 437126 507654 437160
rect 507710 437126 507744 437160
rect 507800 437126 507834 437160
rect 507890 437126 507924 437160
rect 507980 437126 508014 437160
rect 508070 437126 508104 437160
rect 508160 437126 508194 437160
rect 508250 437126 508284 437160
rect 508340 437126 508374 437160
rect 508430 437126 508464 437160
rect 508638 437126 508672 437160
rect 508728 437126 508762 437160
rect 508818 437126 508852 437160
rect 508908 437126 508942 437160
rect 508998 437126 509032 437160
rect 509088 437126 509122 437160
rect 509178 437126 509212 437160
rect 509268 437126 509302 437160
rect 509358 437126 509392 437160
rect 509448 437126 509482 437160
rect 509538 437126 509572 437160
rect 509628 437126 509662 437160
rect 509718 437126 509752 437160
rect 509926 437126 509960 437160
rect 510016 437126 510050 437160
rect 510106 437126 510140 437160
rect 510196 437126 510230 437160
rect 510286 437126 510320 437160
rect 510376 437126 510410 437160
rect 510466 437126 510500 437160
rect 510556 437126 510590 437160
rect 510646 437126 510680 437160
rect 510736 437126 510770 437160
rect 510826 437126 510860 437160
rect 510916 437126 510950 437160
rect 511006 437126 511040 437160
rect 511214 437126 511248 437160
rect 511304 437126 511338 437160
rect 511394 437126 511428 437160
rect 511484 437126 511518 437160
rect 511574 437126 511608 437160
rect 511664 437126 511698 437160
rect 511754 437126 511788 437160
rect 511844 437126 511878 437160
rect 511934 437126 511968 437160
rect 512024 437126 512058 437160
rect 512114 437126 512148 437160
rect 512204 437126 512238 437160
rect 512294 437126 512328 437160
rect 512502 437126 512536 437160
rect 512592 437126 512626 437160
rect 512682 437126 512716 437160
rect 512772 437126 512806 437160
rect 512862 437126 512896 437160
rect 512952 437126 512986 437160
rect 513042 437126 513076 437160
rect 513132 437126 513166 437160
rect 513222 437126 513256 437160
rect 513312 437126 513346 437160
rect 513402 437126 513436 437160
rect 513492 437126 513526 437160
rect 513582 437126 513616 437160
rect 503402 437030 503436 437064
rect 503402 436940 503436 436974
rect 503402 436850 503436 436884
rect 503402 436760 503436 436794
rect 503402 436670 503436 436704
rect 503402 436580 503436 436614
rect 503402 436490 503436 436524
rect 503402 436400 503436 436434
rect 503402 436310 503436 436344
rect 503402 436220 503436 436254
rect 503402 436130 503436 436164
rect 503402 436040 503436 436074
rect 504589 437030 504623 437064
rect 504690 437030 504724 437064
rect 504589 436940 504623 436974
rect 504690 436940 504724 436974
rect 504589 436850 504623 436884
rect 504690 436850 504724 436884
rect 504589 436760 504623 436794
rect 504690 436760 504724 436794
rect 504589 436670 504623 436704
rect 504690 436670 504724 436704
rect 504589 436580 504623 436614
rect 504690 436580 504724 436614
rect 504589 436490 504623 436524
rect 504690 436490 504724 436524
rect 504589 436400 504623 436434
rect 504690 436400 504724 436434
rect 504589 436310 504623 436344
rect 504690 436310 504724 436344
rect 504589 436220 504623 436254
rect 504690 436220 504724 436254
rect 504589 436130 504623 436164
rect 504690 436130 504724 436164
rect 504589 436040 504623 436074
rect 504690 436040 504724 436074
rect 505877 437030 505911 437064
rect 505978 437030 506012 437064
rect 505877 436940 505911 436974
rect 505978 436940 506012 436974
rect 505877 436850 505911 436884
rect 505978 436850 506012 436884
rect 505877 436760 505911 436794
rect 505978 436760 506012 436794
rect 505877 436670 505911 436704
rect 505978 436670 506012 436704
rect 505877 436580 505911 436614
rect 505978 436580 506012 436614
rect 505877 436490 505911 436524
rect 505978 436490 506012 436524
rect 505877 436400 505911 436434
rect 505978 436400 506012 436434
rect 505877 436310 505911 436344
rect 505978 436310 506012 436344
rect 505877 436220 505911 436254
rect 505978 436220 506012 436254
rect 505877 436130 505911 436164
rect 505978 436130 506012 436164
rect 505877 436040 505911 436074
rect 505978 436040 506012 436074
rect 507165 437030 507199 437064
rect 507266 437030 507300 437064
rect 507165 436940 507199 436974
rect 507266 436940 507300 436974
rect 507165 436850 507199 436884
rect 507266 436850 507300 436884
rect 507165 436760 507199 436794
rect 507266 436760 507300 436794
rect 507165 436670 507199 436704
rect 507266 436670 507300 436704
rect 507165 436580 507199 436614
rect 507266 436580 507300 436614
rect 507165 436490 507199 436524
rect 507266 436490 507300 436524
rect 507165 436400 507199 436434
rect 507266 436400 507300 436434
rect 507165 436310 507199 436344
rect 507266 436310 507300 436344
rect 507165 436220 507199 436254
rect 507266 436220 507300 436254
rect 507165 436130 507199 436164
rect 507266 436130 507300 436164
rect 507165 436040 507199 436074
rect 507266 436040 507300 436074
rect 508453 437030 508487 437064
rect 508554 437030 508588 437064
rect 508453 436940 508487 436974
rect 508554 436940 508588 436974
rect 508453 436850 508487 436884
rect 508554 436850 508588 436884
rect 508453 436760 508487 436794
rect 508554 436760 508588 436794
rect 508453 436670 508487 436704
rect 508554 436670 508588 436704
rect 508453 436580 508487 436614
rect 508554 436580 508588 436614
rect 508453 436490 508487 436524
rect 508554 436490 508588 436524
rect 508453 436400 508487 436434
rect 508554 436400 508588 436434
rect 508453 436310 508487 436344
rect 508554 436310 508588 436344
rect 508453 436220 508487 436254
rect 508554 436220 508588 436254
rect 508453 436130 508487 436164
rect 508554 436130 508588 436164
rect 508453 436040 508487 436074
rect 508554 436040 508588 436074
rect 509741 437030 509775 437064
rect 509842 437030 509876 437064
rect 509741 436940 509775 436974
rect 509842 436940 509876 436974
rect 509741 436850 509775 436884
rect 509842 436850 509876 436884
rect 509741 436760 509775 436794
rect 509842 436760 509876 436794
rect 509741 436670 509775 436704
rect 509842 436670 509876 436704
rect 509741 436580 509775 436614
rect 509842 436580 509876 436614
rect 509741 436490 509775 436524
rect 509842 436490 509876 436524
rect 509741 436400 509775 436434
rect 509842 436400 509876 436434
rect 509741 436310 509775 436344
rect 509842 436310 509876 436344
rect 509741 436220 509775 436254
rect 509842 436220 509876 436254
rect 509741 436130 509775 436164
rect 509842 436130 509876 436164
rect 509741 436040 509775 436074
rect 509842 436040 509876 436074
rect 511029 437030 511063 437064
rect 511130 437030 511164 437064
rect 511029 436940 511063 436974
rect 511130 436940 511164 436974
rect 511029 436850 511063 436884
rect 511130 436850 511164 436884
rect 511029 436760 511063 436794
rect 511130 436760 511164 436794
rect 511029 436670 511063 436704
rect 511130 436670 511164 436704
rect 511029 436580 511063 436614
rect 511130 436580 511164 436614
rect 511029 436490 511063 436524
rect 511130 436490 511164 436524
rect 511029 436400 511063 436434
rect 511130 436400 511164 436434
rect 511029 436310 511063 436344
rect 511130 436310 511164 436344
rect 511029 436220 511063 436254
rect 511130 436220 511164 436254
rect 511029 436130 511063 436164
rect 511130 436130 511164 436164
rect 511029 436040 511063 436074
rect 511130 436040 511164 436074
rect 512317 437030 512351 437064
rect 512418 437030 512452 437064
rect 512317 436940 512351 436974
rect 512418 436940 512452 436974
rect 512317 436850 512351 436884
rect 512418 436850 512452 436884
rect 512317 436760 512351 436794
rect 512418 436760 512452 436794
rect 512317 436670 512351 436704
rect 512418 436670 512452 436704
rect 512317 436580 512351 436614
rect 512418 436580 512452 436614
rect 512317 436490 512351 436524
rect 512418 436490 512452 436524
rect 512317 436400 512351 436434
rect 512418 436400 512452 436434
rect 512317 436310 512351 436344
rect 512418 436310 512452 436344
rect 512317 436220 512351 436254
rect 512418 436220 512452 436254
rect 512317 436130 512351 436164
rect 512418 436130 512452 436164
rect 512317 436040 512351 436074
rect 512418 436040 512452 436074
rect 513605 437030 513639 437064
rect 513605 436940 513639 436974
rect 513605 436850 513639 436884
rect 513605 436760 513639 436794
rect 513605 436670 513639 436704
rect 513605 436580 513639 436614
rect 513605 436490 513639 436524
rect 513605 436400 513639 436434
rect 513605 436310 513639 436344
rect 513605 436220 513639 436254
rect 513605 436130 513639 436164
rect 513605 436040 513639 436074
rect 503486 435939 503520 435973
rect 503576 435939 503610 435973
rect 503666 435939 503700 435973
rect 503756 435939 503790 435973
rect 503846 435939 503880 435973
rect 503936 435939 503970 435973
rect 504026 435939 504060 435973
rect 504116 435939 504150 435973
rect 504206 435939 504240 435973
rect 504296 435939 504330 435973
rect 504386 435939 504420 435973
rect 504476 435939 504510 435973
rect 504566 435939 504600 435973
rect 504774 435939 504808 435973
rect 504864 435939 504898 435973
rect 504954 435939 504988 435973
rect 505044 435939 505078 435973
rect 505134 435939 505168 435973
rect 505224 435939 505258 435973
rect 505314 435939 505348 435973
rect 505404 435939 505438 435973
rect 505494 435939 505528 435973
rect 505584 435939 505618 435973
rect 505674 435939 505708 435973
rect 505764 435939 505798 435973
rect 505854 435939 505888 435973
rect 506062 435939 506096 435973
rect 506152 435939 506186 435973
rect 506242 435939 506276 435973
rect 506332 435939 506366 435973
rect 506422 435939 506456 435973
rect 506512 435939 506546 435973
rect 506602 435939 506636 435973
rect 506692 435939 506726 435973
rect 506782 435939 506816 435973
rect 506872 435939 506906 435973
rect 506962 435939 506996 435973
rect 507052 435939 507086 435973
rect 507142 435939 507176 435973
rect 507350 435939 507384 435973
rect 507440 435939 507474 435973
rect 507530 435939 507564 435973
rect 507620 435939 507654 435973
rect 507710 435939 507744 435973
rect 507800 435939 507834 435973
rect 507890 435939 507924 435973
rect 507980 435939 508014 435973
rect 508070 435939 508104 435973
rect 508160 435939 508194 435973
rect 508250 435939 508284 435973
rect 508340 435939 508374 435973
rect 508430 435939 508464 435973
rect 508638 435939 508672 435973
rect 508728 435939 508762 435973
rect 508818 435939 508852 435973
rect 508908 435939 508942 435973
rect 508998 435939 509032 435973
rect 509088 435939 509122 435973
rect 509178 435939 509212 435973
rect 509268 435939 509302 435973
rect 509358 435939 509392 435973
rect 509448 435939 509482 435973
rect 509538 435939 509572 435973
rect 509628 435939 509662 435973
rect 509718 435939 509752 435973
rect 509926 435939 509960 435973
rect 510016 435939 510050 435973
rect 510106 435939 510140 435973
rect 510196 435939 510230 435973
rect 510286 435939 510320 435973
rect 510376 435939 510410 435973
rect 510466 435939 510500 435973
rect 510556 435939 510590 435973
rect 510646 435939 510680 435973
rect 510736 435939 510770 435973
rect 510826 435939 510860 435973
rect 510916 435939 510950 435973
rect 511006 435939 511040 435973
rect 511214 435939 511248 435973
rect 511304 435939 511338 435973
rect 511394 435939 511428 435973
rect 511484 435939 511518 435973
rect 511574 435939 511608 435973
rect 511664 435939 511698 435973
rect 511754 435939 511788 435973
rect 511844 435939 511878 435973
rect 511934 435939 511968 435973
rect 512024 435939 512058 435973
rect 512114 435939 512148 435973
rect 512204 435939 512238 435973
rect 512294 435939 512328 435973
rect 512502 435939 512536 435973
rect 512592 435939 512626 435973
rect 512682 435939 512716 435973
rect 512772 435939 512806 435973
rect 512862 435939 512896 435973
rect 512952 435939 512986 435973
rect 513042 435939 513076 435973
rect 513132 435939 513166 435973
rect 513222 435939 513256 435973
rect 513312 435939 513346 435973
rect 513402 435939 513436 435973
rect 513492 435939 513526 435973
rect 513582 435939 513616 435973
rect 503486 435838 503520 435872
rect 503576 435838 503610 435872
rect 503666 435838 503700 435872
rect 503756 435838 503790 435872
rect 503846 435838 503880 435872
rect 503936 435838 503970 435872
rect 504026 435838 504060 435872
rect 504116 435838 504150 435872
rect 504206 435838 504240 435872
rect 504296 435838 504330 435872
rect 504386 435838 504420 435872
rect 504476 435838 504510 435872
rect 504566 435838 504600 435872
rect 504774 435838 504808 435872
rect 504864 435838 504898 435872
rect 504954 435838 504988 435872
rect 505044 435838 505078 435872
rect 505134 435838 505168 435872
rect 505224 435838 505258 435872
rect 505314 435838 505348 435872
rect 505404 435838 505438 435872
rect 505494 435838 505528 435872
rect 505584 435838 505618 435872
rect 505674 435838 505708 435872
rect 505764 435838 505798 435872
rect 505854 435838 505888 435872
rect 506062 435838 506096 435872
rect 506152 435838 506186 435872
rect 506242 435838 506276 435872
rect 506332 435838 506366 435872
rect 506422 435838 506456 435872
rect 506512 435838 506546 435872
rect 506602 435838 506636 435872
rect 506692 435838 506726 435872
rect 506782 435838 506816 435872
rect 506872 435838 506906 435872
rect 506962 435838 506996 435872
rect 507052 435838 507086 435872
rect 507142 435838 507176 435872
rect 507350 435838 507384 435872
rect 507440 435838 507474 435872
rect 507530 435838 507564 435872
rect 507620 435838 507654 435872
rect 507710 435838 507744 435872
rect 507800 435838 507834 435872
rect 507890 435838 507924 435872
rect 507980 435838 508014 435872
rect 508070 435838 508104 435872
rect 508160 435838 508194 435872
rect 508250 435838 508284 435872
rect 508340 435838 508374 435872
rect 508430 435838 508464 435872
rect 508638 435838 508672 435872
rect 508728 435838 508762 435872
rect 508818 435838 508852 435872
rect 508908 435838 508942 435872
rect 508998 435838 509032 435872
rect 509088 435838 509122 435872
rect 509178 435838 509212 435872
rect 509268 435838 509302 435872
rect 509358 435838 509392 435872
rect 509448 435838 509482 435872
rect 509538 435838 509572 435872
rect 509628 435838 509662 435872
rect 509718 435838 509752 435872
rect 509926 435838 509960 435872
rect 510016 435838 510050 435872
rect 510106 435838 510140 435872
rect 510196 435838 510230 435872
rect 510286 435838 510320 435872
rect 510376 435838 510410 435872
rect 510466 435838 510500 435872
rect 510556 435838 510590 435872
rect 510646 435838 510680 435872
rect 510736 435838 510770 435872
rect 510826 435838 510860 435872
rect 510916 435838 510950 435872
rect 511006 435838 511040 435872
rect 511214 435838 511248 435872
rect 511304 435838 511338 435872
rect 511394 435838 511428 435872
rect 511484 435838 511518 435872
rect 511574 435838 511608 435872
rect 511664 435838 511698 435872
rect 511754 435838 511788 435872
rect 511844 435838 511878 435872
rect 511934 435838 511968 435872
rect 512024 435838 512058 435872
rect 512114 435838 512148 435872
rect 512204 435838 512238 435872
rect 512294 435838 512328 435872
rect 512502 435838 512536 435872
rect 512592 435838 512626 435872
rect 512682 435838 512716 435872
rect 512772 435838 512806 435872
rect 512862 435838 512896 435872
rect 512952 435838 512986 435872
rect 513042 435838 513076 435872
rect 513132 435838 513166 435872
rect 513222 435838 513256 435872
rect 513312 435838 513346 435872
rect 513402 435838 513436 435872
rect 513492 435838 513526 435872
rect 513582 435838 513616 435872
rect 503402 435742 503436 435776
rect 503402 435652 503436 435686
rect 503402 435562 503436 435596
rect 503402 435472 503436 435506
rect 503402 435382 503436 435416
rect 503402 435292 503436 435326
rect 503402 435202 503436 435236
rect 503402 435112 503436 435146
rect 503402 435022 503436 435056
rect 503402 434932 503436 434966
rect 503402 434842 503436 434876
rect 503402 434752 503436 434786
rect 504589 435742 504623 435776
rect 504690 435742 504724 435776
rect 504589 435652 504623 435686
rect 504690 435652 504724 435686
rect 504589 435562 504623 435596
rect 504690 435562 504724 435596
rect 504589 435472 504623 435506
rect 504690 435472 504724 435506
rect 504589 435382 504623 435416
rect 504690 435382 504724 435416
rect 504589 435292 504623 435326
rect 504690 435292 504724 435326
rect 504589 435202 504623 435236
rect 504690 435202 504724 435236
rect 504589 435112 504623 435146
rect 504690 435112 504724 435146
rect 504589 435022 504623 435056
rect 504690 435022 504724 435056
rect 504589 434932 504623 434966
rect 504690 434932 504724 434966
rect 504589 434842 504623 434876
rect 504690 434842 504724 434876
rect 504589 434752 504623 434786
rect 504690 434752 504724 434786
rect 505877 435742 505911 435776
rect 505978 435742 506012 435776
rect 505877 435652 505911 435686
rect 505978 435652 506012 435686
rect 505877 435562 505911 435596
rect 505978 435562 506012 435596
rect 505877 435472 505911 435506
rect 505978 435472 506012 435506
rect 505877 435382 505911 435416
rect 505978 435382 506012 435416
rect 505877 435292 505911 435326
rect 505978 435292 506012 435326
rect 505877 435202 505911 435236
rect 505978 435202 506012 435236
rect 505877 435112 505911 435146
rect 505978 435112 506012 435146
rect 505877 435022 505911 435056
rect 505978 435022 506012 435056
rect 505877 434932 505911 434966
rect 505978 434932 506012 434966
rect 505877 434842 505911 434876
rect 505978 434842 506012 434876
rect 505877 434752 505911 434786
rect 505978 434752 506012 434786
rect 507165 435742 507199 435776
rect 507266 435742 507300 435776
rect 507165 435652 507199 435686
rect 507266 435652 507300 435686
rect 507165 435562 507199 435596
rect 507266 435562 507300 435596
rect 507165 435472 507199 435506
rect 507266 435472 507300 435506
rect 507165 435382 507199 435416
rect 507266 435382 507300 435416
rect 507165 435292 507199 435326
rect 507266 435292 507300 435326
rect 507165 435202 507199 435236
rect 507266 435202 507300 435236
rect 507165 435112 507199 435146
rect 507266 435112 507300 435146
rect 507165 435022 507199 435056
rect 507266 435022 507300 435056
rect 507165 434932 507199 434966
rect 507266 434932 507300 434966
rect 507165 434842 507199 434876
rect 507266 434842 507300 434876
rect 507165 434752 507199 434786
rect 507266 434752 507300 434786
rect 508453 435742 508487 435776
rect 508554 435742 508588 435776
rect 508453 435652 508487 435686
rect 508554 435652 508588 435686
rect 508453 435562 508487 435596
rect 508554 435562 508588 435596
rect 508453 435472 508487 435506
rect 508554 435472 508588 435506
rect 508453 435382 508487 435416
rect 508554 435382 508588 435416
rect 508453 435292 508487 435326
rect 508554 435292 508588 435326
rect 508453 435202 508487 435236
rect 508554 435202 508588 435236
rect 508453 435112 508487 435146
rect 508554 435112 508588 435146
rect 508453 435022 508487 435056
rect 508554 435022 508588 435056
rect 508453 434932 508487 434966
rect 508554 434932 508588 434966
rect 508453 434842 508487 434876
rect 508554 434842 508588 434876
rect 508453 434752 508487 434786
rect 508554 434752 508588 434786
rect 509741 435742 509775 435776
rect 509842 435742 509876 435776
rect 509741 435652 509775 435686
rect 509842 435652 509876 435686
rect 509741 435562 509775 435596
rect 509842 435562 509876 435596
rect 509741 435472 509775 435506
rect 509842 435472 509876 435506
rect 509741 435382 509775 435416
rect 509842 435382 509876 435416
rect 509741 435292 509775 435326
rect 509842 435292 509876 435326
rect 509741 435202 509775 435236
rect 509842 435202 509876 435236
rect 509741 435112 509775 435146
rect 509842 435112 509876 435146
rect 509741 435022 509775 435056
rect 509842 435022 509876 435056
rect 509741 434932 509775 434966
rect 509842 434932 509876 434966
rect 509741 434842 509775 434876
rect 509842 434842 509876 434876
rect 509741 434752 509775 434786
rect 509842 434752 509876 434786
rect 511029 435742 511063 435776
rect 511130 435742 511164 435776
rect 511029 435652 511063 435686
rect 511130 435652 511164 435686
rect 511029 435562 511063 435596
rect 511130 435562 511164 435596
rect 511029 435472 511063 435506
rect 511130 435472 511164 435506
rect 511029 435382 511063 435416
rect 511130 435382 511164 435416
rect 511029 435292 511063 435326
rect 511130 435292 511164 435326
rect 511029 435202 511063 435236
rect 511130 435202 511164 435236
rect 511029 435112 511063 435146
rect 511130 435112 511164 435146
rect 511029 435022 511063 435056
rect 511130 435022 511164 435056
rect 511029 434932 511063 434966
rect 511130 434932 511164 434966
rect 511029 434842 511063 434876
rect 511130 434842 511164 434876
rect 511029 434752 511063 434786
rect 511130 434752 511164 434786
rect 512317 435742 512351 435776
rect 512418 435742 512452 435776
rect 512317 435652 512351 435686
rect 512418 435652 512452 435686
rect 512317 435562 512351 435596
rect 512418 435562 512452 435596
rect 512317 435472 512351 435506
rect 512418 435472 512452 435506
rect 512317 435382 512351 435416
rect 512418 435382 512452 435416
rect 512317 435292 512351 435326
rect 512418 435292 512452 435326
rect 512317 435202 512351 435236
rect 512418 435202 512452 435236
rect 512317 435112 512351 435146
rect 512418 435112 512452 435146
rect 512317 435022 512351 435056
rect 512418 435022 512452 435056
rect 512317 434932 512351 434966
rect 512418 434932 512452 434966
rect 512317 434842 512351 434876
rect 512418 434842 512452 434876
rect 512317 434752 512351 434786
rect 512418 434752 512452 434786
rect 513605 435742 513639 435776
rect 513605 435652 513639 435686
rect 513605 435562 513639 435596
rect 513605 435472 513639 435506
rect 513605 435382 513639 435416
rect 513605 435292 513639 435326
rect 513605 435202 513639 435236
rect 513605 435112 513639 435146
rect 513605 435022 513639 435056
rect 513605 434932 513639 434966
rect 513605 434842 513639 434876
rect 513605 434752 513639 434786
rect 503486 434651 503520 434685
rect 503576 434651 503610 434685
rect 503666 434651 503700 434685
rect 503756 434651 503790 434685
rect 503846 434651 503880 434685
rect 503936 434651 503970 434685
rect 504026 434651 504060 434685
rect 504116 434651 504150 434685
rect 504206 434651 504240 434685
rect 504296 434651 504330 434685
rect 504386 434651 504420 434685
rect 504476 434651 504510 434685
rect 504566 434651 504600 434685
rect 504774 434651 504808 434685
rect 504864 434651 504898 434685
rect 504954 434651 504988 434685
rect 505044 434651 505078 434685
rect 505134 434651 505168 434685
rect 505224 434651 505258 434685
rect 505314 434651 505348 434685
rect 505404 434651 505438 434685
rect 505494 434651 505528 434685
rect 505584 434651 505618 434685
rect 505674 434651 505708 434685
rect 505764 434651 505798 434685
rect 505854 434651 505888 434685
rect 506062 434651 506096 434685
rect 506152 434651 506186 434685
rect 506242 434651 506276 434685
rect 506332 434651 506366 434685
rect 506422 434651 506456 434685
rect 506512 434651 506546 434685
rect 506602 434651 506636 434685
rect 506692 434651 506726 434685
rect 506782 434651 506816 434685
rect 506872 434651 506906 434685
rect 506962 434651 506996 434685
rect 507052 434651 507086 434685
rect 507142 434651 507176 434685
rect 507350 434651 507384 434685
rect 507440 434651 507474 434685
rect 507530 434651 507564 434685
rect 507620 434651 507654 434685
rect 507710 434651 507744 434685
rect 507800 434651 507834 434685
rect 507890 434651 507924 434685
rect 507980 434651 508014 434685
rect 508070 434651 508104 434685
rect 508160 434651 508194 434685
rect 508250 434651 508284 434685
rect 508340 434651 508374 434685
rect 508430 434651 508464 434685
rect 508638 434651 508672 434685
rect 508728 434651 508762 434685
rect 508818 434651 508852 434685
rect 508908 434651 508942 434685
rect 508998 434651 509032 434685
rect 509088 434651 509122 434685
rect 509178 434651 509212 434685
rect 509268 434651 509302 434685
rect 509358 434651 509392 434685
rect 509448 434651 509482 434685
rect 509538 434651 509572 434685
rect 509628 434651 509662 434685
rect 509718 434651 509752 434685
rect 509926 434651 509960 434685
rect 510016 434651 510050 434685
rect 510106 434651 510140 434685
rect 510196 434651 510230 434685
rect 510286 434651 510320 434685
rect 510376 434651 510410 434685
rect 510466 434651 510500 434685
rect 510556 434651 510590 434685
rect 510646 434651 510680 434685
rect 510736 434651 510770 434685
rect 510826 434651 510860 434685
rect 510916 434651 510950 434685
rect 511006 434651 511040 434685
rect 511214 434651 511248 434685
rect 511304 434651 511338 434685
rect 511394 434651 511428 434685
rect 511484 434651 511518 434685
rect 511574 434651 511608 434685
rect 511664 434651 511698 434685
rect 511754 434651 511788 434685
rect 511844 434651 511878 434685
rect 511934 434651 511968 434685
rect 512024 434651 512058 434685
rect 512114 434651 512148 434685
rect 512204 434651 512238 434685
rect 512294 434651 512328 434685
rect 512502 434651 512536 434685
rect 512592 434651 512626 434685
rect 512682 434651 512716 434685
rect 512772 434651 512806 434685
rect 512862 434651 512896 434685
rect 512952 434651 512986 434685
rect 513042 434651 513076 434685
rect 513132 434651 513166 434685
rect 513222 434651 513256 434685
rect 513312 434651 513346 434685
rect 513402 434651 513436 434685
rect 513492 434651 513526 434685
rect 513582 434651 513616 434685
rect 503486 434550 503520 434584
rect 503576 434550 503610 434584
rect 503666 434550 503700 434584
rect 503756 434550 503790 434584
rect 503846 434550 503880 434584
rect 503936 434550 503970 434584
rect 504026 434550 504060 434584
rect 504116 434550 504150 434584
rect 504206 434550 504240 434584
rect 504296 434550 504330 434584
rect 504386 434550 504420 434584
rect 504476 434550 504510 434584
rect 504566 434550 504600 434584
rect 504774 434550 504808 434584
rect 504864 434550 504898 434584
rect 504954 434550 504988 434584
rect 505044 434550 505078 434584
rect 505134 434550 505168 434584
rect 505224 434550 505258 434584
rect 505314 434550 505348 434584
rect 505404 434550 505438 434584
rect 505494 434550 505528 434584
rect 505584 434550 505618 434584
rect 505674 434550 505708 434584
rect 505764 434550 505798 434584
rect 505854 434550 505888 434584
rect 506062 434550 506096 434584
rect 506152 434550 506186 434584
rect 506242 434550 506276 434584
rect 506332 434550 506366 434584
rect 506422 434550 506456 434584
rect 506512 434550 506546 434584
rect 506602 434550 506636 434584
rect 506692 434550 506726 434584
rect 506782 434550 506816 434584
rect 506872 434550 506906 434584
rect 506962 434550 506996 434584
rect 507052 434550 507086 434584
rect 507142 434550 507176 434584
rect 507350 434550 507384 434584
rect 507440 434550 507474 434584
rect 507530 434550 507564 434584
rect 507620 434550 507654 434584
rect 507710 434550 507744 434584
rect 507800 434550 507834 434584
rect 507890 434550 507924 434584
rect 507980 434550 508014 434584
rect 508070 434550 508104 434584
rect 508160 434550 508194 434584
rect 508250 434550 508284 434584
rect 508340 434550 508374 434584
rect 508430 434550 508464 434584
rect 508638 434550 508672 434584
rect 508728 434550 508762 434584
rect 508818 434550 508852 434584
rect 508908 434550 508942 434584
rect 508998 434550 509032 434584
rect 509088 434550 509122 434584
rect 509178 434550 509212 434584
rect 509268 434550 509302 434584
rect 509358 434550 509392 434584
rect 509448 434550 509482 434584
rect 509538 434550 509572 434584
rect 509628 434550 509662 434584
rect 509718 434550 509752 434584
rect 509926 434550 509960 434584
rect 510016 434550 510050 434584
rect 510106 434550 510140 434584
rect 510196 434550 510230 434584
rect 510286 434550 510320 434584
rect 510376 434550 510410 434584
rect 510466 434550 510500 434584
rect 510556 434550 510590 434584
rect 510646 434550 510680 434584
rect 510736 434550 510770 434584
rect 510826 434550 510860 434584
rect 510916 434550 510950 434584
rect 511006 434550 511040 434584
rect 511214 434550 511248 434584
rect 511304 434550 511338 434584
rect 511394 434550 511428 434584
rect 511484 434550 511518 434584
rect 511574 434550 511608 434584
rect 511664 434550 511698 434584
rect 511754 434550 511788 434584
rect 511844 434550 511878 434584
rect 511934 434550 511968 434584
rect 512024 434550 512058 434584
rect 512114 434550 512148 434584
rect 512204 434550 512238 434584
rect 512294 434550 512328 434584
rect 512502 434550 512536 434584
rect 512592 434550 512626 434584
rect 512682 434550 512716 434584
rect 512772 434550 512806 434584
rect 512862 434550 512896 434584
rect 512952 434550 512986 434584
rect 513042 434550 513076 434584
rect 513132 434550 513166 434584
rect 513222 434550 513256 434584
rect 513312 434550 513346 434584
rect 513402 434550 513436 434584
rect 513492 434550 513526 434584
rect 513582 434550 513616 434584
rect 503402 434454 503436 434488
rect 503402 434364 503436 434398
rect 503402 434274 503436 434308
rect 503402 434184 503436 434218
rect 503402 434094 503436 434128
rect 503402 434004 503436 434038
rect 503402 433914 503436 433948
rect 503402 433824 503436 433858
rect 503402 433734 503436 433768
rect 503402 433644 503436 433678
rect 503402 433554 503436 433588
rect 503402 433464 503436 433498
rect 504589 434454 504623 434488
rect 504690 434454 504724 434488
rect 504589 434364 504623 434398
rect 504690 434364 504724 434398
rect 504589 434274 504623 434308
rect 504690 434274 504724 434308
rect 504589 434184 504623 434218
rect 504690 434184 504724 434218
rect 504589 434094 504623 434128
rect 504690 434094 504724 434128
rect 504589 434004 504623 434038
rect 504690 434004 504724 434038
rect 504589 433914 504623 433948
rect 504690 433914 504724 433948
rect 504589 433824 504623 433858
rect 504690 433824 504724 433858
rect 504589 433734 504623 433768
rect 504690 433734 504724 433768
rect 504589 433644 504623 433678
rect 504690 433644 504724 433678
rect 504589 433554 504623 433588
rect 504690 433554 504724 433588
rect 504589 433464 504623 433498
rect 504690 433464 504724 433498
rect 505877 434454 505911 434488
rect 505978 434454 506012 434488
rect 505877 434364 505911 434398
rect 505978 434364 506012 434398
rect 505877 434274 505911 434308
rect 505978 434274 506012 434308
rect 505877 434184 505911 434218
rect 505978 434184 506012 434218
rect 505877 434094 505911 434128
rect 505978 434094 506012 434128
rect 505877 434004 505911 434038
rect 505978 434004 506012 434038
rect 505877 433914 505911 433948
rect 505978 433914 506012 433948
rect 505877 433824 505911 433858
rect 505978 433824 506012 433858
rect 505877 433734 505911 433768
rect 505978 433734 506012 433768
rect 505877 433644 505911 433678
rect 505978 433644 506012 433678
rect 505877 433554 505911 433588
rect 505978 433554 506012 433588
rect 505877 433464 505911 433498
rect 505978 433464 506012 433498
rect 507165 434454 507199 434488
rect 507266 434454 507300 434488
rect 507165 434364 507199 434398
rect 507266 434364 507300 434398
rect 507165 434274 507199 434308
rect 507266 434274 507300 434308
rect 507165 434184 507199 434218
rect 507266 434184 507300 434218
rect 507165 434094 507199 434128
rect 507266 434094 507300 434128
rect 507165 434004 507199 434038
rect 507266 434004 507300 434038
rect 507165 433914 507199 433948
rect 507266 433914 507300 433948
rect 507165 433824 507199 433858
rect 507266 433824 507300 433858
rect 507165 433734 507199 433768
rect 507266 433734 507300 433768
rect 507165 433644 507199 433678
rect 507266 433644 507300 433678
rect 507165 433554 507199 433588
rect 507266 433554 507300 433588
rect 507165 433464 507199 433498
rect 507266 433464 507300 433498
rect 508453 434454 508487 434488
rect 508554 434454 508588 434488
rect 508453 434364 508487 434398
rect 508554 434364 508588 434398
rect 508453 434274 508487 434308
rect 508554 434274 508588 434308
rect 508453 434184 508487 434218
rect 508554 434184 508588 434218
rect 508453 434094 508487 434128
rect 508554 434094 508588 434128
rect 508453 434004 508487 434038
rect 508554 434004 508588 434038
rect 508453 433914 508487 433948
rect 508554 433914 508588 433948
rect 508453 433824 508487 433858
rect 508554 433824 508588 433858
rect 508453 433734 508487 433768
rect 508554 433734 508588 433768
rect 508453 433644 508487 433678
rect 508554 433644 508588 433678
rect 508453 433554 508487 433588
rect 508554 433554 508588 433588
rect 508453 433464 508487 433498
rect 508554 433464 508588 433498
rect 509741 434454 509775 434488
rect 509842 434454 509876 434488
rect 509741 434364 509775 434398
rect 509842 434364 509876 434398
rect 509741 434274 509775 434308
rect 509842 434274 509876 434308
rect 509741 434184 509775 434218
rect 509842 434184 509876 434218
rect 509741 434094 509775 434128
rect 509842 434094 509876 434128
rect 509741 434004 509775 434038
rect 509842 434004 509876 434038
rect 509741 433914 509775 433948
rect 509842 433914 509876 433948
rect 509741 433824 509775 433858
rect 509842 433824 509876 433858
rect 509741 433734 509775 433768
rect 509842 433734 509876 433768
rect 509741 433644 509775 433678
rect 509842 433644 509876 433678
rect 509741 433554 509775 433588
rect 509842 433554 509876 433588
rect 509741 433464 509775 433498
rect 509842 433464 509876 433498
rect 511029 434454 511063 434488
rect 511130 434454 511164 434488
rect 511029 434364 511063 434398
rect 511130 434364 511164 434398
rect 511029 434274 511063 434308
rect 511130 434274 511164 434308
rect 511029 434184 511063 434218
rect 511130 434184 511164 434218
rect 511029 434094 511063 434128
rect 511130 434094 511164 434128
rect 511029 434004 511063 434038
rect 511130 434004 511164 434038
rect 511029 433914 511063 433948
rect 511130 433914 511164 433948
rect 511029 433824 511063 433858
rect 511130 433824 511164 433858
rect 511029 433734 511063 433768
rect 511130 433734 511164 433768
rect 511029 433644 511063 433678
rect 511130 433644 511164 433678
rect 511029 433554 511063 433588
rect 511130 433554 511164 433588
rect 511029 433464 511063 433498
rect 511130 433464 511164 433498
rect 512317 434454 512351 434488
rect 512418 434454 512452 434488
rect 512317 434364 512351 434398
rect 512418 434364 512452 434398
rect 512317 434274 512351 434308
rect 512418 434274 512452 434308
rect 512317 434184 512351 434218
rect 512418 434184 512452 434218
rect 512317 434094 512351 434128
rect 512418 434094 512452 434128
rect 512317 434004 512351 434038
rect 512418 434004 512452 434038
rect 512317 433914 512351 433948
rect 512418 433914 512452 433948
rect 512317 433824 512351 433858
rect 512418 433824 512452 433858
rect 512317 433734 512351 433768
rect 512418 433734 512452 433768
rect 512317 433644 512351 433678
rect 512418 433644 512452 433678
rect 512317 433554 512351 433588
rect 512418 433554 512452 433588
rect 512317 433464 512351 433498
rect 512418 433464 512452 433498
rect 513605 434454 513639 434488
rect 513605 434364 513639 434398
rect 513605 434274 513639 434308
rect 513605 434184 513639 434218
rect 513605 434094 513639 434128
rect 513605 434004 513639 434038
rect 513605 433914 513639 433948
rect 513605 433824 513639 433858
rect 513605 433734 513639 433768
rect 513605 433644 513639 433678
rect 513605 433554 513639 433588
rect 513605 433464 513639 433498
rect 503486 433363 503520 433397
rect 503576 433363 503610 433397
rect 503666 433363 503700 433397
rect 503756 433363 503790 433397
rect 503846 433363 503880 433397
rect 503936 433363 503970 433397
rect 504026 433363 504060 433397
rect 504116 433363 504150 433397
rect 504206 433363 504240 433397
rect 504296 433363 504330 433397
rect 504386 433363 504420 433397
rect 504476 433363 504510 433397
rect 504566 433363 504600 433397
rect 504774 433363 504808 433397
rect 504864 433363 504898 433397
rect 504954 433363 504988 433397
rect 505044 433363 505078 433397
rect 505134 433363 505168 433397
rect 505224 433363 505258 433397
rect 505314 433363 505348 433397
rect 505404 433363 505438 433397
rect 505494 433363 505528 433397
rect 505584 433363 505618 433397
rect 505674 433363 505708 433397
rect 505764 433363 505798 433397
rect 505854 433363 505888 433397
rect 506062 433363 506096 433397
rect 506152 433363 506186 433397
rect 506242 433363 506276 433397
rect 506332 433363 506366 433397
rect 506422 433363 506456 433397
rect 506512 433363 506546 433397
rect 506602 433363 506636 433397
rect 506692 433363 506726 433397
rect 506782 433363 506816 433397
rect 506872 433363 506906 433397
rect 506962 433363 506996 433397
rect 507052 433363 507086 433397
rect 507142 433363 507176 433397
rect 507350 433363 507384 433397
rect 507440 433363 507474 433397
rect 507530 433363 507564 433397
rect 507620 433363 507654 433397
rect 507710 433363 507744 433397
rect 507800 433363 507834 433397
rect 507890 433363 507924 433397
rect 507980 433363 508014 433397
rect 508070 433363 508104 433397
rect 508160 433363 508194 433397
rect 508250 433363 508284 433397
rect 508340 433363 508374 433397
rect 508430 433363 508464 433397
rect 508638 433363 508672 433397
rect 508728 433363 508762 433397
rect 508818 433363 508852 433397
rect 508908 433363 508942 433397
rect 508998 433363 509032 433397
rect 509088 433363 509122 433397
rect 509178 433363 509212 433397
rect 509268 433363 509302 433397
rect 509358 433363 509392 433397
rect 509448 433363 509482 433397
rect 509538 433363 509572 433397
rect 509628 433363 509662 433397
rect 509718 433363 509752 433397
rect 509926 433363 509960 433397
rect 510016 433363 510050 433397
rect 510106 433363 510140 433397
rect 510196 433363 510230 433397
rect 510286 433363 510320 433397
rect 510376 433363 510410 433397
rect 510466 433363 510500 433397
rect 510556 433363 510590 433397
rect 510646 433363 510680 433397
rect 510736 433363 510770 433397
rect 510826 433363 510860 433397
rect 510916 433363 510950 433397
rect 511006 433363 511040 433397
rect 511214 433363 511248 433397
rect 511304 433363 511338 433397
rect 511394 433363 511428 433397
rect 511484 433363 511518 433397
rect 511574 433363 511608 433397
rect 511664 433363 511698 433397
rect 511754 433363 511788 433397
rect 511844 433363 511878 433397
rect 511934 433363 511968 433397
rect 512024 433363 512058 433397
rect 512114 433363 512148 433397
rect 512204 433363 512238 433397
rect 512294 433363 512328 433397
rect 512502 433363 512536 433397
rect 512592 433363 512626 433397
rect 512682 433363 512716 433397
rect 512772 433363 512806 433397
rect 512862 433363 512896 433397
rect 512952 433363 512986 433397
rect 513042 433363 513076 433397
rect 513132 433363 513166 433397
rect 513222 433363 513256 433397
rect 513312 433363 513346 433397
rect 513402 433363 513436 433397
rect 513492 433363 513526 433397
rect 513582 433363 513616 433397
rect 503486 433262 503520 433296
rect 503576 433262 503610 433296
rect 503666 433262 503700 433296
rect 503756 433262 503790 433296
rect 503846 433262 503880 433296
rect 503936 433262 503970 433296
rect 504026 433262 504060 433296
rect 504116 433262 504150 433296
rect 504206 433262 504240 433296
rect 504296 433262 504330 433296
rect 504386 433262 504420 433296
rect 504476 433262 504510 433296
rect 504566 433262 504600 433296
rect 504774 433262 504808 433296
rect 504864 433262 504898 433296
rect 504954 433262 504988 433296
rect 505044 433262 505078 433296
rect 505134 433262 505168 433296
rect 505224 433262 505258 433296
rect 505314 433262 505348 433296
rect 505404 433262 505438 433296
rect 505494 433262 505528 433296
rect 505584 433262 505618 433296
rect 505674 433262 505708 433296
rect 505764 433262 505798 433296
rect 505854 433262 505888 433296
rect 506062 433262 506096 433296
rect 506152 433262 506186 433296
rect 506242 433262 506276 433296
rect 506332 433262 506366 433296
rect 506422 433262 506456 433296
rect 506512 433262 506546 433296
rect 506602 433262 506636 433296
rect 506692 433262 506726 433296
rect 506782 433262 506816 433296
rect 506872 433262 506906 433296
rect 506962 433262 506996 433296
rect 507052 433262 507086 433296
rect 507142 433262 507176 433296
rect 507350 433262 507384 433296
rect 507440 433262 507474 433296
rect 507530 433262 507564 433296
rect 507620 433262 507654 433296
rect 507710 433262 507744 433296
rect 507800 433262 507834 433296
rect 507890 433262 507924 433296
rect 507980 433262 508014 433296
rect 508070 433262 508104 433296
rect 508160 433262 508194 433296
rect 508250 433262 508284 433296
rect 508340 433262 508374 433296
rect 508430 433262 508464 433296
rect 508638 433262 508672 433296
rect 508728 433262 508762 433296
rect 508818 433262 508852 433296
rect 508908 433262 508942 433296
rect 508998 433262 509032 433296
rect 509088 433262 509122 433296
rect 509178 433262 509212 433296
rect 509268 433262 509302 433296
rect 509358 433262 509392 433296
rect 509448 433262 509482 433296
rect 509538 433262 509572 433296
rect 509628 433262 509662 433296
rect 509718 433262 509752 433296
rect 509926 433262 509960 433296
rect 510016 433262 510050 433296
rect 510106 433262 510140 433296
rect 510196 433262 510230 433296
rect 510286 433262 510320 433296
rect 510376 433262 510410 433296
rect 510466 433262 510500 433296
rect 510556 433262 510590 433296
rect 510646 433262 510680 433296
rect 510736 433262 510770 433296
rect 510826 433262 510860 433296
rect 510916 433262 510950 433296
rect 511006 433262 511040 433296
rect 511214 433262 511248 433296
rect 511304 433262 511338 433296
rect 511394 433262 511428 433296
rect 511484 433262 511518 433296
rect 511574 433262 511608 433296
rect 511664 433262 511698 433296
rect 511754 433262 511788 433296
rect 511844 433262 511878 433296
rect 511934 433262 511968 433296
rect 512024 433262 512058 433296
rect 512114 433262 512148 433296
rect 512204 433262 512238 433296
rect 512294 433262 512328 433296
rect 512502 433262 512536 433296
rect 512592 433262 512626 433296
rect 512682 433262 512716 433296
rect 512772 433262 512806 433296
rect 512862 433262 512896 433296
rect 512952 433262 512986 433296
rect 513042 433262 513076 433296
rect 513132 433262 513166 433296
rect 513222 433262 513256 433296
rect 513312 433262 513346 433296
rect 513402 433262 513436 433296
rect 513492 433262 513526 433296
rect 513582 433262 513616 433296
rect 503402 433166 503436 433200
rect 503402 433076 503436 433110
rect 503402 432986 503436 433020
rect 503402 432896 503436 432930
rect 503402 432806 503436 432840
rect 503402 432716 503436 432750
rect 503402 432626 503436 432660
rect 503402 432536 503436 432570
rect 503402 432446 503436 432480
rect 503402 432356 503436 432390
rect 503402 432266 503436 432300
rect 503402 432176 503436 432210
rect 504589 433166 504623 433200
rect 504690 433166 504724 433200
rect 504589 433076 504623 433110
rect 504690 433076 504724 433110
rect 504589 432986 504623 433020
rect 504690 432986 504724 433020
rect 504589 432896 504623 432930
rect 504690 432896 504724 432930
rect 504589 432806 504623 432840
rect 504690 432806 504724 432840
rect 504589 432716 504623 432750
rect 504690 432716 504724 432750
rect 504589 432626 504623 432660
rect 504690 432626 504724 432660
rect 504589 432536 504623 432570
rect 504690 432536 504724 432570
rect 504589 432446 504623 432480
rect 504690 432446 504724 432480
rect 504589 432356 504623 432390
rect 504690 432356 504724 432390
rect 504589 432266 504623 432300
rect 504690 432266 504724 432300
rect 504589 432176 504623 432210
rect 504690 432176 504724 432210
rect 505877 433166 505911 433200
rect 505978 433166 506012 433200
rect 505877 433076 505911 433110
rect 505978 433076 506012 433110
rect 505877 432986 505911 433020
rect 505978 432986 506012 433020
rect 505877 432896 505911 432930
rect 505978 432896 506012 432930
rect 505877 432806 505911 432840
rect 505978 432806 506012 432840
rect 505877 432716 505911 432750
rect 505978 432716 506012 432750
rect 505877 432626 505911 432660
rect 505978 432626 506012 432660
rect 505877 432536 505911 432570
rect 505978 432536 506012 432570
rect 505877 432446 505911 432480
rect 505978 432446 506012 432480
rect 505877 432356 505911 432390
rect 505978 432356 506012 432390
rect 505877 432266 505911 432300
rect 505978 432266 506012 432300
rect 505877 432176 505911 432210
rect 505978 432176 506012 432210
rect 507165 433166 507199 433200
rect 507266 433166 507300 433200
rect 507165 433076 507199 433110
rect 507266 433076 507300 433110
rect 507165 432986 507199 433020
rect 507266 432986 507300 433020
rect 507165 432896 507199 432930
rect 507266 432896 507300 432930
rect 507165 432806 507199 432840
rect 507266 432806 507300 432840
rect 507165 432716 507199 432750
rect 507266 432716 507300 432750
rect 507165 432626 507199 432660
rect 507266 432626 507300 432660
rect 507165 432536 507199 432570
rect 507266 432536 507300 432570
rect 507165 432446 507199 432480
rect 507266 432446 507300 432480
rect 507165 432356 507199 432390
rect 507266 432356 507300 432390
rect 507165 432266 507199 432300
rect 507266 432266 507300 432300
rect 507165 432176 507199 432210
rect 507266 432176 507300 432210
rect 508453 433166 508487 433200
rect 508554 433166 508588 433200
rect 508453 433076 508487 433110
rect 508554 433076 508588 433110
rect 508453 432986 508487 433020
rect 508554 432986 508588 433020
rect 508453 432896 508487 432930
rect 508554 432896 508588 432930
rect 508453 432806 508487 432840
rect 508554 432806 508588 432840
rect 508453 432716 508487 432750
rect 508554 432716 508588 432750
rect 508453 432626 508487 432660
rect 508554 432626 508588 432660
rect 508453 432536 508487 432570
rect 508554 432536 508588 432570
rect 508453 432446 508487 432480
rect 508554 432446 508588 432480
rect 508453 432356 508487 432390
rect 508554 432356 508588 432390
rect 508453 432266 508487 432300
rect 508554 432266 508588 432300
rect 508453 432176 508487 432210
rect 508554 432176 508588 432210
rect 509741 433166 509775 433200
rect 509842 433166 509876 433200
rect 509741 433076 509775 433110
rect 509842 433076 509876 433110
rect 509741 432986 509775 433020
rect 509842 432986 509876 433020
rect 509741 432896 509775 432930
rect 509842 432896 509876 432930
rect 509741 432806 509775 432840
rect 509842 432806 509876 432840
rect 509741 432716 509775 432750
rect 509842 432716 509876 432750
rect 509741 432626 509775 432660
rect 509842 432626 509876 432660
rect 509741 432536 509775 432570
rect 509842 432536 509876 432570
rect 509741 432446 509775 432480
rect 509842 432446 509876 432480
rect 509741 432356 509775 432390
rect 509842 432356 509876 432390
rect 509741 432266 509775 432300
rect 509842 432266 509876 432300
rect 509741 432176 509775 432210
rect 509842 432176 509876 432210
rect 511029 433166 511063 433200
rect 511130 433166 511164 433200
rect 511029 433076 511063 433110
rect 511130 433076 511164 433110
rect 511029 432986 511063 433020
rect 511130 432986 511164 433020
rect 511029 432896 511063 432930
rect 511130 432896 511164 432930
rect 511029 432806 511063 432840
rect 511130 432806 511164 432840
rect 511029 432716 511063 432750
rect 511130 432716 511164 432750
rect 511029 432626 511063 432660
rect 511130 432626 511164 432660
rect 511029 432536 511063 432570
rect 511130 432536 511164 432570
rect 511029 432446 511063 432480
rect 511130 432446 511164 432480
rect 511029 432356 511063 432390
rect 511130 432356 511164 432390
rect 511029 432266 511063 432300
rect 511130 432266 511164 432300
rect 511029 432176 511063 432210
rect 511130 432176 511164 432210
rect 512317 433166 512351 433200
rect 512418 433166 512452 433200
rect 512317 433076 512351 433110
rect 512418 433076 512452 433110
rect 512317 432986 512351 433020
rect 512418 432986 512452 433020
rect 512317 432896 512351 432930
rect 512418 432896 512452 432930
rect 512317 432806 512351 432840
rect 512418 432806 512452 432840
rect 512317 432716 512351 432750
rect 512418 432716 512452 432750
rect 512317 432626 512351 432660
rect 512418 432626 512452 432660
rect 512317 432536 512351 432570
rect 512418 432536 512452 432570
rect 512317 432446 512351 432480
rect 512418 432446 512452 432480
rect 512317 432356 512351 432390
rect 512418 432356 512452 432390
rect 512317 432266 512351 432300
rect 512418 432266 512452 432300
rect 512317 432176 512351 432210
rect 512418 432176 512452 432210
rect 513605 433166 513639 433200
rect 513605 433076 513639 433110
rect 513605 432986 513639 433020
rect 513605 432896 513639 432930
rect 513605 432806 513639 432840
rect 513605 432716 513639 432750
rect 513605 432626 513639 432660
rect 513605 432536 513639 432570
rect 513605 432446 513639 432480
rect 513605 432356 513639 432390
rect 513605 432266 513639 432300
rect 513605 432176 513639 432210
rect 503486 432075 503520 432109
rect 503576 432075 503610 432109
rect 503666 432075 503700 432109
rect 503756 432075 503790 432109
rect 503846 432075 503880 432109
rect 503936 432075 503970 432109
rect 504026 432075 504060 432109
rect 504116 432075 504150 432109
rect 504206 432075 504240 432109
rect 504296 432075 504330 432109
rect 504386 432075 504420 432109
rect 504476 432075 504510 432109
rect 504566 432075 504600 432109
rect 504774 432075 504808 432109
rect 504864 432075 504898 432109
rect 504954 432075 504988 432109
rect 505044 432075 505078 432109
rect 505134 432075 505168 432109
rect 505224 432075 505258 432109
rect 505314 432075 505348 432109
rect 505404 432075 505438 432109
rect 505494 432075 505528 432109
rect 505584 432075 505618 432109
rect 505674 432075 505708 432109
rect 505764 432075 505798 432109
rect 505854 432075 505888 432109
rect 506062 432075 506096 432109
rect 506152 432075 506186 432109
rect 506242 432075 506276 432109
rect 506332 432075 506366 432109
rect 506422 432075 506456 432109
rect 506512 432075 506546 432109
rect 506602 432075 506636 432109
rect 506692 432075 506726 432109
rect 506782 432075 506816 432109
rect 506872 432075 506906 432109
rect 506962 432075 506996 432109
rect 507052 432075 507086 432109
rect 507142 432075 507176 432109
rect 507350 432075 507384 432109
rect 507440 432075 507474 432109
rect 507530 432075 507564 432109
rect 507620 432075 507654 432109
rect 507710 432075 507744 432109
rect 507800 432075 507834 432109
rect 507890 432075 507924 432109
rect 507980 432075 508014 432109
rect 508070 432075 508104 432109
rect 508160 432075 508194 432109
rect 508250 432075 508284 432109
rect 508340 432075 508374 432109
rect 508430 432075 508464 432109
rect 508638 432075 508672 432109
rect 508728 432075 508762 432109
rect 508818 432075 508852 432109
rect 508908 432075 508942 432109
rect 508998 432075 509032 432109
rect 509088 432075 509122 432109
rect 509178 432075 509212 432109
rect 509268 432075 509302 432109
rect 509358 432075 509392 432109
rect 509448 432075 509482 432109
rect 509538 432075 509572 432109
rect 509628 432075 509662 432109
rect 509718 432075 509752 432109
rect 509926 432075 509960 432109
rect 510016 432075 510050 432109
rect 510106 432075 510140 432109
rect 510196 432075 510230 432109
rect 510286 432075 510320 432109
rect 510376 432075 510410 432109
rect 510466 432075 510500 432109
rect 510556 432075 510590 432109
rect 510646 432075 510680 432109
rect 510736 432075 510770 432109
rect 510826 432075 510860 432109
rect 510916 432075 510950 432109
rect 511006 432075 511040 432109
rect 511214 432075 511248 432109
rect 511304 432075 511338 432109
rect 511394 432075 511428 432109
rect 511484 432075 511518 432109
rect 511574 432075 511608 432109
rect 511664 432075 511698 432109
rect 511754 432075 511788 432109
rect 511844 432075 511878 432109
rect 511934 432075 511968 432109
rect 512024 432075 512058 432109
rect 512114 432075 512148 432109
rect 512204 432075 512238 432109
rect 512294 432075 512328 432109
rect 512502 432075 512536 432109
rect 512592 432075 512626 432109
rect 512682 432075 512716 432109
rect 512772 432075 512806 432109
rect 512862 432075 512896 432109
rect 512952 432075 512986 432109
rect 513042 432075 513076 432109
rect 513132 432075 513166 432109
rect 513222 432075 513256 432109
rect 513312 432075 513346 432109
rect 513402 432075 513436 432109
rect 513492 432075 513526 432109
rect 513582 432075 513616 432109
rect 500344 430044 526568 431044
rect 527592 430020 528592 475332
rect 572412 455212 577642 455246
rect 572316 454056 572350 455150
rect 577704 454056 577738 455150
rect 572412 453960 577642 453994
<< nsubdiffcont >>
rect 562252 495480 567482 495514
rect 562156 494315 562190 495417
rect 567544 494315 567578 495417
rect 562252 494218 567482 494252
rect 503226 470102 505568 470202
rect 502622 464278 502722 466620
rect 503226 460974 505568 461074
rect 503528 460052 510528 460252
rect 503528 454142 510528 454342
rect 503528 448642 510528 448842
rect 503526 442686 510526 442886
rect 503665 438266 503699 438300
rect 503755 438266 503789 438300
rect 503845 438266 503879 438300
rect 503935 438266 503969 438300
rect 504025 438266 504059 438300
rect 504115 438266 504149 438300
rect 504205 438266 504239 438300
rect 504295 438266 504329 438300
rect 504385 438266 504419 438300
rect 503552 438188 503586 438222
rect 503552 438098 503586 438132
rect 503552 438008 503586 438042
rect 503552 437918 503586 437952
rect 503552 437828 503586 437862
rect 503552 437738 503586 437772
rect 503552 437648 503586 437682
rect 503552 437558 503586 437592
rect 503552 437468 503586 437502
rect 504442 438154 504476 438188
rect 504442 438064 504476 438098
rect 504442 437974 504476 438008
rect 504442 437884 504476 437918
rect 504442 437794 504476 437828
rect 504442 437704 504476 437738
rect 504442 437614 504476 437648
rect 504442 437524 504476 437558
rect 504442 437434 504476 437468
rect 503646 437376 503680 437410
rect 503736 437376 503770 437410
rect 503826 437376 503860 437410
rect 503916 437376 503950 437410
rect 504006 437376 504040 437410
rect 504096 437376 504130 437410
rect 504186 437376 504220 437410
rect 504276 437376 504310 437410
rect 504366 437376 504400 437410
rect 504953 438266 504987 438300
rect 505043 438266 505077 438300
rect 505133 438266 505167 438300
rect 505223 438266 505257 438300
rect 505313 438266 505347 438300
rect 505403 438266 505437 438300
rect 505493 438266 505527 438300
rect 505583 438266 505617 438300
rect 505673 438266 505707 438300
rect 504840 438188 504874 438222
rect 504840 438098 504874 438132
rect 504840 438008 504874 438042
rect 504840 437918 504874 437952
rect 504840 437828 504874 437862
rect 504840 437738 504874 437772
rect 504840 437648 504874 437682
rect 504840 437558 504874 437592
rect 504840 437468 504874 437502
rect 505730 438154 505764 438188
rect 505730 438064 505764 438098
rect 505730 437974 505764 438008
rect 505730 437884 505764 437918
rect 505730 437794 505764 437828
rect 505730 437704 505764 437738
rect 505730 437614 505764 437648
rect 505730 437524 505764 437558
rect 505730 437434 505764 437468
rect 504934 437376 504968 437410
rect 505024 437376 505058 437410
rect 505114 437376 505148 437410
rect 505204 437376 505238 437410
rect 505294 437376 505328 437410
rect 505384 437376 505418 437410
rect 505474 437376 505508 437410
rect 505564 437376 505598 437410
rect 505654 437376 505688 437410
rect 506241 438266 506275 438300
rect 506331 438266 506365 438300
rect 506421 438266 506455 438300
rect 506511 438266 506545 438300
rect 506601 438266 506635 438300
rect 506691 438266 506725 438300
rect 506781 438266 506815 438300
rect 506871 438266 506905 438300
rect 506961 438266 506995 438300
rect 506128 438188 506162 438222
rect 506128 438098 506162 438132
rect 506128 438008 506162 438042
rect 506128 437918 506162 437952
rect 506128 437828 506162 437862
rect 506128 437738 506162 437772
rect 506128 437648 506162 437682
rect 506128 437558 506162 437592
rect 506128 437468 506162 437502
rect 507018 438154 507052 438188
rect 507018 438064 507052 438098
rect 507018 437974 507052 438008
rect 507018 437884 507052 437918
rect 507018 437794 507052 437828
rect 507018 437704 507052 437738
rect 507018 437614 507052 437648
rect 507018 437524 507052 437558
rect 507018 437434 507052 437468
rect 506222 437376 506256 437410
rect 506312 437376 506346 437410
rect 506402 437376 506436 437410
rect 506492 437376 506526 437410
rect 506582 437376 506616 437410
rect 506672 437376 506706 437410
rect 506762 437376 506796 437410
rect 506852 437376 506886 437410
rect 506942 437376 506976 437410
rect 507529 438266 507563 438300
rect 507619 438266 507653 438300
rect 507709 438266 507743 438300
rect 507799 438266 507833 438300
rect 507889 438266 507923 438300
rect 507979 438266 508013 438300
rect 508069 438266 508103 438300
rect 508159 438266 508193 438300
rect 508249 438266 508283 438300
rect 507416 438188 507450 438222
rect 507416 438098 507450 438132
rect 507416 438008 507450 438042
rect 507416 437918 507450 437952
rect 507416 437828 507450 437862
rect 507416 437738 507450 437772
rect 507416 437648 507450 437682
rect 507416 437558 507450 437592
rect 507416 437468 507450 437502
rect 508306 438154 508340 438188
rect 508306 438064 508340 438098
rect 508306 437974 508340 438008
rect 508306 437884 508340 437918
rect 508306 437794 508340 437828
rect 508306 437704 508340 437738
rect 508306 437614 508340 437648
rect 508306 437524 508340 437558
rect 508306 437434 508340 437468
rect 507510 437376 507544 437410
rect 507600 437376 507634 437410
rect 507690 437376 507724 437410
rect 507780 437376 507814 437410
rect 507870 437376 507904 437410
rect 507960 437376 507994 437410
rect 508050 437376 508084 437410
rect 508140 437376 508174 437410
rect 508230 437376 508264 437410
rect 508817 438266 508851 438300
rect 508907 438266 508941 438300
rect 508997 438266 509031 438300
rect 509087 438266 509121 438300
rect 509177 438266 509211 438300
rect 509267 438266 509301 438300
rect 509357 438266 509391 438300
rect 509447 438266 509481 438300
rect 509537 438266 509571 438300
rect 508704 438188 508738 438222
rect 508704 438098 508738 438132
rect 508704 438008 508738 438042
rect 508704 437918 508738 437952
rect 508704 437828 508738 437862
rect 508704 437738 508738 437772
rect 508704 437648 508738 437682
rect 508704 437558 508738 437592
rect 508704 437468 508738 437502
rect 509594 438154 509628 438188
rect 509594 438064 509628 438098
rect 509594 437974 509628 438008
rect 509594 437884 509628 437918
rect 509594 437794 509628 437828
rect 509594 437704 509628 437738
rect 509594 437614 509628 437648
rect 509594 437524 509628 437558
rect 509594 437434 509628 437468
rect 508798 437376 508832 437410
rect 508888 437376 508922 437410
rect 508978 437376 509012 437410
rect 509068 437376 509102 437410
rect 509158 437376 509192 437410
rect 509248 437376 509282 437410
rect 509338 437376 509372 437410
rect 509428 437376 509462 437410
rect 509518 437376 509552 437410
rect 510105 438266 510139 438300
rect 510195 438266 510229 438300
rect 510285 438266 510319 438300
rect 510375 438266 510409 438300
rect 510465 438266 510499 438300
rect 510555 438266 510589 438300
rect 510645 438266 510679 438300
rect 510735 438266 510769 438300
rect 510825 438266 510859 438300
rect 509992 438188 510026 438222
rect 509992 438098 510026 438132
rect 509992 438008 510026 438042
rect 509992 437918 510026 437952
rect 509992 437828 510026 437862
rect 509992 437738 510026 437772
rect 509992 437648 510026 437682
rect 509992 437558 510026 437592
rect 509992 437468 510026 437502
rect 510882 438154 510916 438188
rect 510882 438064 510916 438098
rect 510882 437974 510916 438008
rect 510882 437884 510916 437918
rect 510882 437794 510916 437828
rect 510882 437704 510916 437738
rect 510882 437614 510916 437648
rect 510882 437524 510916 437558
rect 510882 437434 510916 437468
rect 510086 437376 510120 437410
rect 510176 437376 510210 437410
rect 510266 437376 510300 437410
rect 510356 437376 510390 437410
rect 510446 437376 510480 437410
rect 510536 437376 510570 437410
rect 510626 437376 510660 437410
rect 510716 437376 510750 437410
rect 510806 437376 510840 437410
rect 511393 438266 511427 438300
rect 511483 438266 511517 438300
rect 511573 438266 511607 438300
rect 511663 438266 511697 438300
rect 511753 438266 511787 438300
rect 511843 438266 511877 438300
rect 511933 438266 511967 438300
rect 512023 438266 512057 438300
rect 512113 438266 512147 438300
rect 511280 438188 511314 438222
rect 511280 438098 511314 438132
rect 511280 438008 511314 438042
rect 511280 437918 511314 437952
rect 511280 437828 511314 437862
rect 511280 437738 511314 437772
rect 511280 437648 511314 437682
rect 511280 437558 511314 437592
rect 511280 437468 511314 437502
rect 512170 438154 512204 438188
rect 512170 438064 512204 438098
rect 512170 437974 512204 438008
rect 512170 437884 512204 437918
rect 512170 437794 512204 437828
rect 512170 437704 512204 437738
rect 512170 437614 512204 437648
rect 512170 437524 512204 437558
rect 512170 437434 512204 437468
rect 511374 437376 511408 437410
rect 511464 437376 511498 437410
rect 511554 437376 511588 437410
rect 511644 437376 511678 437410
rect 511734 437376 511768 437410
rect 511824 437376 511858 437410
rect 511914 437376 511948 437410
rect 512004 437376 512038 437410
rect 512094 437376 512128 437410
rect 512681 438266 512715 438300
rect 512771 438266 512805 438300
rect 512861 438266 512895 438300
rect 512951 438266 512985 438300
rect 513041 438266 513075 438300
rect 513131 438266 513165 438300
rect 513221 438266 513255 438300
rect 513311 438266 513345 438300
rect 513401 438266 513435 438300
rect 512568 438188 512602 438222
rect 512568 438098 512602 438132
rect 512568 438008 512602 438042
rect 512568 437918 512602 437952
rect 512568 437828 512602 437862
rect 512568 437738 512602 437772
rect 512568 437648 512602 437682
rect 512568 437558 512602 437592
rect 512568 437468 512602 437502
rect 513458 438154 513492 438188
rect 513458 438064 513492 438098
rect 513458 437974 513492 438008
rect 513458 437884 513492 437918
rect 513458 437794 513492 437828
rect 513458 437704 513492 437738
rect 513458 437614 513492 437648
rect 513458 437524 513492 437558
rect 513458 437434 513492 437468
rect 512662 437376 512696 437410
rect 512752 437376 512786 437410
rect 512842 437376 512876 437410
rect 512932 437376 512966 437410
rect 513022 437376 513056 437410
rect 513112 437376 513146 437410
rect 513202 437376 513236 437410
rect 513292 437376 513326 437410
rect 513382 437376 513416 437410
rect 503665 436978 503699 437012
rect 503755 436978 503789 437012
rect 503845 436978 503879 437012
rect 503935 436978 503969 437012
rect 504025 436978 504059 437012
rect 504115 436978 504149 437012
rect 504205 436978 504239 437012
rect 504295 436978 504329 437012
rect 504385 436978 504419 437012
rect 503552 436900 503586 436934
rect 503552 436810 503586 436844
rect 503552 436720 503586 436754
rect 503552 436630 503586 436664
rect 503552 436540 503586 436574
rect 503552 436450 503586 436484
rect 503552 436360 503586 436394
rect 503552 436270 503586 436304
rect 503552 436180 503586 436214
rect 504442 436866 504476 436900
rect 504442 436776 504476 436810
rect 504442 436686 504476 436720
rect 504442 436596 504476 436630
rect 504442 436506 504476 436540
rect 504442 436416 504476 436450
rect 504442 436326 504476 436360
rect 504442 436236 504476 436270
rect 504442 436146 504476 436180
rect 503646 436088 503680 436122
rect 503736 436088 503770 436122
rect 503826 436088 503860 436122
rect 503916 436088 503950 436122
rect 504006 436088 504040 436122
rect 504096 436088 504130 436122
rect 504186 436088 504220 436122
rect 504276 436088 504310 436122
rect 504366 436088 504400 436122
rect 504953 436978 504987 437012
rect 505043 436978 505077 437012
rect 505133 436978 505167 437012
rect 505223 436978 505257 437012
rect 505313 436978 505347 437012
rect 505403 436978 505437 437012
rect 505493 436978 505527 437012
rect 505583 436978 505617 437012
rect 505673 436978 505707 437012
rect 504840 436900 504874 436934
rect 504840 436810 504874 436844
rect 504840 436720 504874 436754
rect 504840 436630 504874 436664
rect 504840 436540 504874 436574
rect 504840 436450 504874 436484
rect 504840 436360 504874 436394
rect 504840 436270 504874 436304
rect 504840 436180 504874 436214
rect 505730 436866 505764 436900
rect 505730 436776 505764 436810
rect 505730 436686 505764 436720
rect 505730 436596 505764 436630
rect 505730 436506 505764 436540
rect 505730 436416 505764 436450
rect 505730 436326 505764 436360
rect 505730 436236 505764 436270
rect 505730 436146 505764 436180
rect 504934 436088 504968 436122
rect 505024 436088 505058 436122
rect 505114 436088 505148 436122
rect 505204 436088 505238 436122
rect 505294 436088 505328 436122
rect 505384 436088 505418 436122
rect 505474 436088 505508 436122
rect 505564 436088 505598 436122
rect 505654 436088 505688 436122
rect 506241 436978 506275 437012
rect 506331 436978 506365 437012
rect 506421 436978 506455 437012
rect 506511 436978 506545 437012
rect 506601 436978 506635 437012
rect 506691 436978 506725 437012
rect 506781 436978 506815 437012
rect 506871 436978 506905 437012
rect 506961 436978 506995 437012
rect 506128 436900 506162 436934
rect 506128 436810 506162 436844
rect 506128 436720 506162 436754
rect 506128 436630 506162 436664
rect 506128 436540 506162 436574
rect 506128 436450 506162 436484
rect 506128 436360 506162 436394
rect 506128 436270 506162 436304
rect 506128 436180 506162 436214
rect 507018 436866 507052 436900
rect 507018 436776 507052 436810
rect 507018 436686 507052 436720
rect 507018 436596 507052 436630
rect 507018 436506 507052 436540
rect 507018 436416 507052 436450
rect 507018 436326 507052 436360
rect 507018 436236 507052 436270
rect 507018 436146 507052 436180
rect 506222 436088 506256 436122
rect 506312 436088 506346 436122
rect 506402 436088 506436 436122
rect 506492 436088 506526 436122
rect 506582 436088 506616 436122
rect 506672 436088 506706 436122
rect 506762 436088 506796 436122
rect 506852 436088 506886 436122
rect 506942 436088 506976 436122
rect 507529 436978 507563 437012
rect 507619 436978 507653 437012
rect 507709 436978 507743 437012
rect 507799 436978 507833 437012
rect 507889 436978 507923 437012
rect 507979 436978 508013 437012
rect 508069 436978 508103 437012
rect 508159 436978 508193 437012
rect 508249 436978 508283 437012
rect 507416 436900 507450 436934
rect 507416 436810 507450 436844
rect 507416 436720 507450 436754
rect 507416 436630 507450 436664
rect 507416 436540 507450 436574
rect 507416 436450 507450 436484
rect 507416 436360 507450 436394
rect 507416 436270 507450 436304
rect 507416 436180 507450 436214
rect 508306 436866 508340 436900
rect 508306 436776 508340 436810
rect 508306 436686 508340 436720
rect 508306 436596 508340 436630
rect 508306 436506 508340 436540
rect 508306 436416 508340 436450
rect 508306 436326 508340 436360
rect 508306 436236 508340 436270
rect 508306 436146 508340 436180
rect 507510 436088 507544 436122
rect 507600 436088 507634 436122
rect 507690 436088 507724 436122
rect 507780 436088 507814 436122
rect 507870 436088 507904 436122
rect 507960 436088 507994 436122
rect 508050 436088 508084 436122
rect 508140 436088 508174 436122
rect 508230 436088 508264 436122
rect 508817 436978 508851 437012
rect 508907 436978 508941 437012
rect 508997 436978 509031 437012
rect 509087 436978 509121 437012
rect 509177 436978 509211 437012
rect 509267 436978 509301 437012
rect 509357 436978 509391 437012
rect 509447 436978 509481 437012
rect 509537 436978 509571 437012
rect 508704 436900 508738 436934
rect 508704 436810 508738 436844
rect 508704 436720 508738 436754
rect 508704 436630 508738 436664
rect 508704 436540 508738 436574
rect 508704 436450 508738 436484
rect 508704 436360 508738 436394
rect 508704 436270 508738 436304
rect 508704 436180 508738 436214
rect 509594 436866 509628 436900
rect 509594 436776 509628 436810
rect 509594 436686 509628 436720
rect 509594 436596 509628 436630
rect 509594 436506 509628 436540
rect 509594 436416 509628 436450
rect 509594 436326 509628 436360
rect 509594 436236 509628 436270
rect 509594 436146 509628 436180
rect 508798 436088 508832 436122
rect 508888 436088 508922 436122
rect 508978 436088 509012 436122
rect 509068 436088 509102 436122
rect 509158 436088 509192 436122
rect 509248 436088 509282 436122
rect 509338 436088 509372 436122
rect 509428 436088 509462 436122
rect 509518 436088 509552 436122
rect 510105 436978 510139 437012
rect 510195 436978 510229 437012
rect 510285 436978 510319 437012
rect 510375 436978 510409 437012
rect 510465 436978 510499 437012
rect 510555 436978 510589 437012
rect 510645 436978 510679 437012
rect 510735 436978 510769 437012
rect 510825 436978 510859 437012
rect 509992 436900 510026 436934
rect 509992 436810 510026 436844
rect 509992 436720 510026 436754
rect 509992 436630 510026 436664
rect 509992 436540 510026 436574
rect 509992 436450 510026 436484
rect 509992 436360 510026 436394
rect 509992 436270 510026 436304
rect 509992 436180 510026 436214
rect 510882 436866 510916 436900
rect 510882 436776 510916 436810
rect 510882 436686 510916 436720
rect 510882 436596 510916 436630
rect 510882 436506 510916 436540
rect 510882 436416 510916 436450
rect 510882 436326 510916 436360
rect 510882 436236 510916 436270
rect 510882 436146 510916 436180
rect 510086 436088 510120 436122
rect 510176 436088 510210 436122
rect 510266 436088 510300 436122
rect 510356 436088 510390 436122
rect 510446 436088 510480 436122
rect 510536 436088 510570 436122
rect 510626 436088 510660 436122
rect 510716 436088 510750 436122
rect 510806 436088 510840 436122
rect 511393 436978 511427 437012
rect 511483 436978 511517 437012
rect 511573 436978 511607 437012
rect 511663 436978 511697 437012
rect 511753 436978 511787 437012
rect 511843 436978 511877 437012
rect 511933 436978 511967 437012
rect 512023 436978 512057 437012
rect 512113 436978 512147 437012
rect 511280 436900 511314 436934
rect 511280 436810 511314 436844
rect 511280 436720 511314 436754
rect 511280 436630 511314 436664
rect 511280 436540 511314 436574
rect 511280 436450 511314 436484
rect 511280 436360 511314 436394
rect 511280 436270 511314 436304
rect 511280 436180 511314 436214
rect 512170 436866 512204 436900
rect 512170 436776 512204 436810
rect 512170 436686 512204 436720
rect 512170 436596 512204 436630
rect 512170 436506 512204 436540
rect 512170 436416 512204 436450
rect 512170 436326 512204 436360
rect 512170 436236 512204 436270
rect 512170 436146 512204 436180
rect 511374 436088 511408 436122
rect 511464 436088 511498 436122
rect 511554 436088 511588 436122
rect 511644 436088 511678 436122
rect 511734 436088 511768 436122
rect 511824 436088 511858 436122
rect 511914 436088 511948 436122
rect 512004 436088 512038 436122
rect 512094 436088 512128 436122
rect 512681 436978 512715 437012
rect 512771 436978 512805 437012
rect 512861 436978 512895 437012
rect 512951 436978 512985 437012
rect 513041 436978 513075 437012
rect 513131 436978 513165 437012
rect 513221 436978 513255 437012
rect 513311 436978 513345 437012
rect 513401 436978 513435 437012
rect 512568 436900 512602 436934
rect 512568 436810 512602 436844
rect 512568 436720 512602 436754
rect 512568 436630 512602 436664
rect 512568 436540 512602 436574
rect 512568 436450 512602 436484
rect 512568 436360 512602 436394
rect 512568 436270 512602 436304
rect 512568 436180 512602 436214
rect 513458 436866 513492 436900
rect 513458 436776 513492 436810
rect 513458 436686 513492 436720
rect 513458 436596 513492 436630
rect 513458 436506 513492 436540
rect 513458 436416 513492 436450
rect 513458 436326 513492 436360
rect 513458 436236 513492 436270
rect 513458 436146 513492 436180
rect 512662 436088 512696 436122
rect 512752 436088 512786 436122
rect 512842 436088 512876 436122
rect 512932 436088 512966 436122
rect 513022 436088 513056 436122
rect 513112 436088 513146 436122
rect 513202 436088 513236 436122
rect 513292 436088 513326 436122
rect 513382 436088 513416 436122
rect 503665 435690 503699 435724
rect 503755 435690 503789 435724
rect 503845 435690 503879 435724
rect 503935 435690 503969 435724
rect 504025 435690 504059 435724
rect 504115 435690 504149 435724
rect 504205 435690 504239 435724
rect 504295 435690 504329 435724
rect 504385 435690 504419 435724
rect 503552 435612 503586 435646
rect 503552 435522 503586 435556
rect 503552 435432 503586 435466
rect 503552 435342 503586 435376
rect 503552 435252 503586 435286
rect 503552 435162 503586 435196
rect 503552 435072 503586 435106
rect 503552 434982 503586 435016
rect 503552 434892 503586 434926
rect 504442 435578 504476 435612
rect 504442 435488 504476 435522
rect 504442 435398 504476 435432
rect 504442 435308 504476 435342
rect 504442 435218 504476 435252
rect 504442 435128 504476 435162
rect 504442 435038 504476 435072
rect 504442 434948 504476 434982
rect 504442 434858 504476 434892
rect 503646 434800 503680 434834
rect 503736 434800 503770 434834
rect 503826 434800 503860 434834
rect 503916 434800 503950 434834
rect 504006 434800 504040 434834
rect 504096 434800 504130 434834
rect 504186 434800 504220 434834
rect 504276 434800 504310 434834
rect 504366 434800 504400 434834
rect 504953 435690 504987 435724
rect 505043 435690 505077 435724
rect 505133 435690 505167 435724
rect 505223 435690 505257 435724
rect 505313 435690 505347 435724
rect 505403 435690 505437 435724
rect 505493 435690 505527 435724
rect 505583 435690 505617 435724
rect 505673 435690 505707 435724
rect 504840 435612 504874 435646
rect 504840 435522 504874 435556
rect 504840 435432 504874 435466
rect 504840 435342 504874 435376
rect 504840 435252 504874 435286
rect 504840 435162 504874 435196
rect 504840 435072 504874 435106
rect 504840 434982 504874 435016
rect 504840 434892 504874 434926
rect 505730 435578 505764 435612
rect 505730 435488 505764 435522
rect 505730 435398 505764 435432
rect 505730 435308 505764 435342
rect 505730 435218 505764 435252
rect 505730 435128 505764 435162
rect 505730 435038 505764 435072
rect 505730 434948 505764 434982
rect 505730 434858 505764 434892
rect 504934 434800 504968 434834
rect 505024 434800 505058 434834
rect 505114 434800 505148 434834
rect 505204 434800 505238 434834
rect 505294 434800 505328 434834
rect 505384 434800 505418 434834
rect 505474 434800 505508 434834
rect 505564 434800 505598 434834
rect 505654 434800 505688 434834
rect 506241 435690 506275 435724
rect 506331 435690 506365 435724
rect 506421 435690 506455 435724
rect 506511 435690 506545 435724
rect 506601 435690 506635 435724
rect 506691 435690 506725 435724
rect 506781 435690 506815 435724
rect 506871 435690 506905 435724
rect 506961 435690 506995 435724
rect 506128 435612 506162 435646
rect 506128 435522 506162 435556
rect 506128 435432 506162 435466
rect 506128 435342 506162 435376
rect 506128 435252 506162 435286
rect 506128 435162 506162 435196
rect 506128 435072 506162 435106
rect 506128 434982 506162 435016
rect 506128 434892 506162 434926
rect 507018 435578 507052 435612
rect 507018 435488 507052 435522
rect 507018 435398 507052 435432
rect 507018 435308 507052 435342
rect 507018 435218 507052 435252
rect 507018 435128 507052 435162
rect 507018 435038 507052 435072
rect 507018 434948 507052 434982
rect 507018 434858 507052 434892
rect 506222 434800 506256 434834
rect 506312 434800 506346 434834
rect 506402 434800 506436 434834
rect 506492 434800 506526 434834
rect 506582 434800 506616 434834
rect 506672 434800 506706 434834
rect 506762 434800 506796 434834
rect 506852 434800 506886 434834
rect 506942 434800 506976 434834
rect 507529 435690 507563 435724
rect 507619 435690 507653 435724
rect 507709 435690 507743 435724
rect 507799 435690 507833 435724
rect 507889 435690 507923 435724
rect 507979 435690 508013 435724
rect 508069 435690 508103 435724
rect 508159 435690 508193 435724
rect 508249 435690 508283 435724
rect 507416 435612 507450 435646
rect 507416 435522 507450 435556
rect 507416 435432 507450 435466
rect 507416 435342 507450 435376
rect 507416 435252 507450 435286
rect 507416 435162 507450 435196
rect 507416 435072 507450 435106
rect 507416 434982 507450 435016
rect 507416 434892 507450 434926
rect 508306 435578 508340 435612
rect 508306 435488 508340 435522
rect 508306 435398 508340 435432
rect 508306 435308 508340 435342
rect 508306 435218 508340 435252
rect 508306 435128 508340 435162
rect 508306 435038 508340 435072
rect 508306 434948 508340 434982
rect 508306 434858 508340 434892
rect 507510 434800 507544 434834
rect 507600 434800 507634 434834
rect 507690 434800 507724 434834
rect 507780 434800 507814 434834
rect 507870 434800 507904 434834
rect 507960 434800 507994 434834
rect 508050 434800 508084 434834
rect 508140 434800 508174 434834
rect 508230 434800 508264 434834
rect 508817 435690 508851 435724
rect 508907 435690 508941 435724
rect 508997 435690 509031 435724
rect 509087 435690 509121 435724
rect 509177 435690 509211 435724
rect 509267 435690 509301 435724
rect 509357 435690 509391 435724
rect 509447 435690 509481 435724
rect 509537 435690 509571 435724
rect 508704 435612 508738 435646
rect 508704 435522 508738 435556
rect 508704 435432 508738 435466
rect 508704 435342 508738 435376
rect 508704 435252 508738 435286
rect 508704 435162 508738 435196
rect 508704 435072 508738 435106
rect 508704 434982 508738 435016
rect 508704 434892 508738 434926
rect 509594 435578 509628 435612
rect 509594 435488 509628 435522
rect 509594 435398 509628 435432
rect 509594 435308 509628 435342
rect 509594 435218 509628 435252
rect 509594 435128 509628 435162
rect 509594 435038 509628 435072
rect 509594 434948 509628 434982
rect 509594 434858 509628 434892
rect 508798 434800 508832 434834
rect 508888 434800 508922 434834
rect 508978 434800 509012 434834
rect 509068 434800 509102 434834
rect 509158 434800 509192 434834
rect 509248 434800 509282 434834
rect 509338 434800 509372 434834
rect 509428 434800 509462 434834
rect 509518 434800 509552 434834
rect 510105 435690 510139 435724
rect 510195 435690 510229 435724
rect 510285 435690 510319 435724
rect 510375 435690 510409 435724
rect 510465 435690 510499 435724
rect 510555 435690 510589 435724
rect 510645 435690 510679 435724
rect 510735 435690 510769 435724
rect 510825 435690 510859 435724
rect 509992 435612 510026 435646
rect 509992 435522 510026 435556
rect 509992 435432 510026 435466
rect 509992 435342 510026 435376
rect 509992 435252 510026 435286
rect 509992 435162 510026 435196
rect 509992 435072 510026 435106
rect 509992 434982 510026 435016
rect 509992 434892 510026 434926
rect 510882 435578 510916 435612
rect 510882 435488 510916 435522
rect 510882 435398 510916 435432
rect 510882 435308 510916 435342
rect 510882 435218 510916 435252
rect 510882 435128 510916 435162
rect 510882 435038 510916 435072
rect 510882 434948 510916 434982
rect 510882 434858 510916 434892
rect 510086 434800 510120 434834
rect 510176 434800 510210 434834
rect 510266 434800 510300 434834
rect 510356 434800 510390 434834
rect 510446 434800 510480 434834
rect 510536 434800 510570 434834
rect 510626 434800 510660 434834
rect 510716 434800 510750 434834
rect 510806 434800 510840 434834
rect 511393 435690 511427 435724
rect 511483 435690 511517 435724
rect 511573 435690 511607 435724
rect 511663 435690 511697 435724
rect 511753 435690 511787 435724
rect 511843 435690 511877 435724
rect 511933 435690 511967 435724
rect 512023 435690 512057 435724
rect 512113 435690 512147 435724
rect 511280 435612 511314 435646
rect 511280 435522 511314 435556
rect 511280 435432 511314 435466
rect 511280 435342 511314 435376
rect 511280 435252 511314 435286
rect 511280 435162 511314 435196
rect 511280 435072 511314 435106
rect 511280 434982 511314 435016
rect 511280 434892 511314 434926
rect 512170 435578 512204 435612
rect 512170 435488 512204 435522
rect 512170 435398 512204 435432
rect 512170 435308 512204 435342
rect 512170 435218 512204 435252
rect 512170 435128 512204 435162
rect 512170 435038 512204 435072
rect 512170 434948 512204 434982
rect 512170 434858 512204 434892
rect 511374 434800 511408 434834
rect 511464 434800 511498 434834
rect 511554 434800 511588 434834
rect 511644 434800 511678 434834
rect 511734 434800 511768 434834
rect 511824 434800 511858 434834
rect 511914 434800 511948 434834
rect 512004 434800 512038 434834
rect 512094 434800 512128 434834
rect 512681 435690 512715 435724
rect 512771 435690 512805 435724
rect 512861 435690 512895 435724
rect 512951 435690 512985 435724
rect 513041 435690 513075 435724
rect 513131 435690 513165 435724
rect 513221 435690 513255 435724
rect 513311 435690 513345 435724
rect 513401 435690 513435 435724
rect 512568 435612 512602 435646
rect 512568 435522 512602 435556
rect 512568 435432 512602 435466
rect 512568 435342 512602 435376
rect 512568 435252 512602 435286
rect 512568 435162 512602 435196
rect 512568 435072 512602 435106
rect 512568 434982 512602 435016
rect 512568 434892 512602 434926
rect 513458 435578 513492 435612
rect 513458 435488 513492 435522
rect 513458 435398 513492 435432
rect 513458 435308 513492 435342
rect 513458 435218 513492 435252
rect 513458 435128 513492 435162
rect 513458 435038 513492 435072
rect 513458 434948 513492 434982
rect 513458 434858 513492 434892
rect 512662 434800 512696 434834
rect 512752 434800 512786 434834
rect 512842 434800 512876 434834
rect 512932 434800 512966 434834
rect 513022 434800 513056 434834
rect 513112 434800 513146 434834
rect 513202 434800 513236 434834
rect 513292 434800 513326 434834
rect 513382 434800 513416 434834
rect 503665 434402 503699 434436
rect 503755 434402 503789 434436
rect 503845 434402 503879 434436
rect 503935 434402 503969 434436
rect 504025 434402 504059 434436
rect 504115 434402 504149 434436
rect 504205 434402 504239 434436
rect 504295 434402 504329 434436
rect 504385 434402 504419 434436
rect 503552 434324 503586 434358
rect 503552 434234 503586 434268
rect 503552 434144 503586 434178
rect 503552 434054 503586 434088
rect 503552 433964 503586 433998
rect 503552 433874 503586 433908
rect 503552 433784 503586 433818
rect 503552 433694 503586 433728
rect 503552 433604 503586 433638
rect 504442 434290 504476 434324
rect 504442 434200 504476 434234
rect 504442 434110 504476 434144
rect 504442 434020 504476 434054
rect 504442 433930 504476 433964
rect 504442 433840 504476 433874
rect 504442 433750 504476 433784
rect 504442 433660 504476 433694
rect 504442 433570 504476 433604
rect 503646 433512 503680 433546
rect 503736 433512 503770 433546
rect 503826 433512 503860 433546
rect 503916 433512 503950 433546
rect 504006 433512 504040 433546
rect 504096 433512 504130 433546
rect 504186 433512 504220 433546
rect 504276 433512 504310 433546
rect 504366 433512 504400 433546
rect 504953 434402 504987 434436
rect 505043 434402 505077 434436
rect 505133 434402 505167 434436
rect 505223 434402 505257 434436
rect 505313 434402 505347 434436
rect 505403 434402 505437 434436
rect 505493 434402 505527 434436
rect 505583 434402 505617 434436
rect 505673 434402 505707 434436
rect 504840 434324 504874 434358
rect 504840 434234 504874 434268
rect 504840 434144 504874 434178
rect 504840 434054 504874 434088
rect 504840 433964 504874 433998
rect 504840 433874 504874 433908
rect 504840 433784 504874 433818
rect 504840 433694 504874 433728
rect 504840 433604 504874 433638
rect 505730 434290 505764 434324
rect 505730 434200 505764 434234
rect 505730 434110 505764 434144
rect 505730 434020 505764 434054
rect 505730 433930 505764 433964
rect 505730 433840 505764 433874
rect 505730 433750 505764 433784
rect 505730 433660 505764 433694
rect 505730 433570 505764 433604
rect 504934 433512 504968 433546
rect 505024 433512 505058 433546
rect 505114 433512 505148 433546
rect 505204 433512 505238 433546
rect 505294 433512 505328 433546
rect 505384 433512 505418 433546
rect 505474 433512 505508 433546
rect 505564 433512 505598 433546
rect 505654 433512 505688 433546
rect 506241 434402 506275 434436
rect 506331 434402 506365 434436
rect 506421 434402 506455 434436
rect 506511 434402 506545 434436
rect 506601 434402 506635 434436
rect 506691 434402 506725 434436
rect 506781 434402 506815 434436
rect 506871 434402 506905 434436
rect 506961 434402 506995 434436
rect 506128 434324 506162 434358
rect 506128 434234 506162 434268
rect 506128 434144 506162 434178
rect 506128 434054 506162 434088
rect 506128 433964 506162 433998
rect 506128 433874 506162 433908
rect 506128 433784 506162 433818
rect 506128 433694 506162 433728
rect 506128 433604 506162 433638
rect 507018 434290 507052 434324
rect 507018 434200 507052 434234
rect 507018 434110 507052 434144
rect 507018 434020 507052 434054
rect 507018 433930 507052 433964
rect 507018 433840 507052 433874
rect 507018 433750 507052 433784
rect 507018 433660 507052 433694
rect 507018 433570 507052 433604
rect 506222 433512 506256 433546
rect 506312 433512 506346 433546
rect 506402 433512 506436 433546
rect 506492 433512 506526 433546
rect 506582 433512 506616 433546
rect 506672 433512 506706 433546
rect 506762 433512 506796 433546
rect 506852 433512 506886 433546
rect 506942 433512 506976 433546
rect 507529 434402 507563 434436
rect 507619 434402 507653 434436
rect 507709 434402 507743 434436
rect 507799 434402 507833 434436
rect 507889 434402 507923 434436
rect 507979 434402 508013 434436
rect 508069 434402 508103 434436
rect 508159 434402 508193 434436
rect 508249 434402 508283 434436
rect 507416 434324 507450 434358
rect 507416 434234 507450 434268
rect 507416 434144 507450 434178
rect 507416 434054 507450 434088
rect 507416 433964 507450 433998
rect 507416 433874 507450 433908
rect 507416 433784 507450 433818
rect 507416 433694 507450 433728
rect 507416 433604 507450 433638
rect 508306 434290 508340 434324
rect 508306 434200 508340 434234
rect 508306 434110 508340 434144
rect 508306 434020 508340 434054
rect 508306 433930 508340 433964
rect 508306 433840 508340 433874
rect 508306 433750 508340 433784
rect 508306 433660 508340 433694
rect 508306 433570 508340 433604
rect 507510 433512 507544 433546
rect 507600 433512 507634 433546
rect 507690 433512 507724 433546
rect 507780 433512 507814 433546
rect 507870 433512 507904 433546
rect 507960 433512 507994 433546
rect 508050 433512 508084 433546
rect 508140 433512 508174 433546
rect 508230 433512 508264 433546
rect 508817 434402 508851 434436
rect 508907 434402 508941 434436
rect 508997 434402 509031 434436
rect 509087 434402 509121 434436
rect 509177 434402 509211 434436
rect 509267 434402 509301 434436
rect 509357 434402 509391 434436
rect 509447 434402 509481 434436
rect 509537 434402 509571 434436
rect 508704 434324 508738 434358
rect 508704 434234 508738 434268
rect 508704 434144 508738 434178
rect 508704 434054 508738 434088
rect 508704 433964 508738 433998
rect 508704 433874 508738 433908
rect 508704 433784 508738 433818
rect 508704 433694 508738 433728
rect 508704 433604 508738 433638
rect 509594 434290 509628 434324
rect 509594 434200 509628 434234
rect 509594 434110 509628 434144
rect 509594 434020 509628 434054
rect 509594 433930 509628 433964
rect 509594 433840 509628 433874
rect 509594 433750 509628 433784
rect 509594 433660 509628 433694
rect 509594 433570 509628 433604
rect 508798 433512 508832 433546
rect 508888 433512 508922 433546
rect 508978 433512 509012 433546
rect 509068 433512 509102 433546
rect 509158 433512 509192 433546
rect 509248 433512 509282 433546
rect 509338 433512 509372 433546
rect 509428 433512 509462 433546
rect 509518 433512 509552 433546
rect 510105 434402 510139 434436
rect 510195 434402 510229 434436
rect 510285 434402 510319 434436
rect 510375 434402 510409 434436
rect 510465 434402 510499 434436
rect 510555 434402 510589 434436
rect 510645 434402 510679 434436
rect 510735 434402 510769 434436
rect 510825 434402 510859 434436
rect 509992 434324 510026 434358
rect 509992 434234 510026 434268
rect 509992 434144 510026 434178
rect 509992 434054 510026 434088
rect 509992 433964 510026 433998
rect 509992 433874 510026 433908
rect 509992 433784 510026 433818
rect 509992 433694 510026 433728
rect 509992 433604 510026 433638
rect 510882 434290 510916 434324
rect 510882 434200 510916 434234
rect 510882 434110 510916 434144
rect 510882 434020 510916 434054
rect 510882 433930 510916 433964
rect 510882 433840 510916 433874
rect 510882 433750 510916 433784
rect 510882 433660 510916 433694
rect 510882 433570 510916 433604
rect 510086 433512 510120 433546
rect 510176 433512 510210 433546
rect 510266 433512 510300 433546
rect 510356 433512 510390 433546
rect 510446 433512 510480 433546
rect 510536 433512 510570 433546
rect 510626 433512 510660 433546
rect 510716 433512 510750 433546
rect 510806 433512 510840 433546
rect 511393 434402 511427 434436
rect 511483 434402 511517 434436
rect 511573 434402 511607 434436
rect 511663 434402 511697 434436
rect 511753 434402 511787 434436
rect 511843 434402 511877 434436
rect 511933 434402 511967 434436
rect 512023 434402 512057 434436
rect 512113 434402 512147 434436
rect 511280 434324 511314 434358
rect 511280 434234 511314 434268
rect 511280 434144 511314 434178
rect 511280 434054 511314 434088
rect 511280 433964 511314 433998
rect 511280 433874 511314 433908
rect 511280 433784 511314 433818
rect 511280 433694 511314 433728
rect 511280 433604 511314 433638
rect 512170 434290 512204 434324
rect 512170 434200 512204 434234
rect 512170 434110 512204 434144
rect 512170 434020 512204 434054
rect 512170 433930 512204 433964
rect 512170 433840 512204 433874
rect 512170 433750 512204 433784
rect 512170 433660 512204 433694
rect 512170 433570 512204 433604
rect 511374 433512 511408 433546
rect 511464 433512 511498 433546
rect 511554 433512 511588 433546
rect 511644 433512 511678 433546
rect 511734 433512 511768 433546
rect 511824 433512 511858 433546
rect 511914 433512 511948 433546
rect 512004 433512 512038 433546
rect 512094 433512 512128 433546
rect 512681 434402 512715 434436
rect 512771 434402 512805 434436
rect 512861 434402 512895 434436
rect 512951 434402 512985 434436
rect 513041 434402 513075 434436
rect 513131 434402 513165 434436
rect 513221 434402 513255 434436
rect 513311 434402 513345 434436
rect 513401 434402 513435 434436
rect 512568 434324 512602 434358
rect 512568 434234 512602 434268
rect 512568 434144 512602 434178
rect 512568 434054 512602 434088
rect 512568 433964 512602 433998
rect 512568 433874 512602 433908
rect 512568 433784 512602 433818
rect 512568 433694 512602 433728
rect 512568 433604 512602 433638
rect 513458 434290 513492 434324
rect 513458 434200 513492 434234
rect 513458 434110 513492 434144
rect 513458 434020 513492 434054
rect 513458 433930 513492 433964
rect 513458 433840 513492 433874
rect 513458 433750 513492 433784
rect 513458 433660 513492 433694
rect 513458 433570 513492 433604
rect 512662 433512 512696 433546
rect 512752 433512 512786 433546
rect 512842 433512 512876 433546
rect 512932 433512 512966 433546
rect 513022 433512 513056 433546
rect 513112 433512 513146 433546
rect 513202 433512 513236 433546
rect 513292 433512 513326 433546
rect 513382 433512 513416 433546
rect 503665 433114 503699 433148
rect 503755 433114 503789 433148
rect 503845 433114 503879 433148
rect 503935 433114 503969 433148
rect 504025 433114 504059 433148
rect 504115 433114 504149 433148
rect 504205 433114 504239 433148
rect 504295 433114 504329 433148
rect 504385 433114 504419 433148
rect 503552 433036 503586 433070
rect 503552 432946 503586 432980
rect 503552 432856 503586 432890
rect 503552 432766 503586 432800
rect 503552 432676 503586 432710
rect 503552 432586 503586 432620
rect 503552 432496 503586 432530
rect 503552 432406 503586 432440
rect 503552 432316 503586 432350
rect 504442 433002 504476 433036
rect 504442 432912 504476 432946
rect 504442 432822 504476 432856
rect 504442 432732 504476 432766
rect 504442 432642 504476 432676
rect 504442 432552 504476 432586
rect 504442 432462 504476 432496
rect 504442 432372 504476 432406
rect 504442 432282 504476 432316
rect 503646 432224 503680 432258
rect 503736 432224 503770 432258
rect 503826 432224 503860 432258
rect 503916 432224 503950 432258
rect 504006 432224 504040 432258
rect 504096 432224 504130 432258
rect 504186 432224 504220 432258
rect 504276 432224 504310 432258
rect 504366 432224 504400 432258
rect 504953 433114 504987 433148
rect 505043 433114 505077 433148
rect 505133 433114 505167 433148
rect 505223 433114 505257 433148
rect 505313 433114 505347 433148
rect 505403 433114 505437 433148
rect 505493 433114 505527 433148
rect 505583 433114 505617 433148
rect 505673 433114 505707 433148
rect 504840 433036 504874 433070
rect 504840 432946 504874 432980
rect 504840 432856 504874 432890
rect 504840 432766 504874 432800
rect 504840 432676 504874 432710
rect 504840 432586 504874 432620
rect 504840 432496 504874 432530
rect 504840 432406 504874 432440
rect 504840 432316 504874 432350
rect 505730 433002 505764 433036
rect 505730 432912 505764 432946
rect 505730 432822 505764 432856
rect 505730 432732 505764 432766
rect 505730 432642 505764 432676
rect 505730 432552 505764 432586
rect 505730 432462 505764 432496
rect 505730 432372 505764 432406
rect 505730 432282 505764 432316
rect 504934 432224 504968 432258
rect 505024 432224 505058 432258
rect 505114 432224 505148 432258
rect 505204 432224 505238 432258
rect 505294 432224 505328 432258
rect 505384 432224 505418 432258
rect 505474 432224 505508 432258
rect 505564 432224 505598 432258
rect 505654 432224 505688 432258
rect 506241 433114 506275 433148
rect 506331 433114 506365 433148
rect 506421 433114 506455 433148
rect 506511 433114 506545 433148
rect 506601 433114 506635 433148
rect 506691 433114 506725 433148
rect 506781 433114 506815 433148
rect 506871 433114 506905 433148
rect 506961 433114 506995 433148
rect 506128 433036 506162 433070
rect 506128 432946 506162 432980
rect 506128 432856 506162 432890
rect 506128 432766 506162 432800
rect 506128 432676 506162 432710
rect 506128 432586 506162 432620
rect 506128 432496 506162 432530
rect 506128 432406 506162 432440
rect 506128 432316 506162 432350
rect 507018 433002 507052 433036
rect 507018 432912 507052 432946
rect 507018 432822 507052 432856
rect 507018 432732 507052 432766
rect 507018 432642 507052 432676
rect 507018 432552 507052 432586
rect 507018 432462 507052 432496
rect 507018 432372 507052 432406
rect 507018 432282 507052 432316
rect 506222 432224 506256 432258
rect 506312 432224 506346 432258
rect 506402 432224 506436 432258
rect 506492 432224 506526 432258
rect 506582 432224 506616 432258
rect 506672 432224 506706 432258
rect 506762 432224 506796 432258
rect 506852 432224 506886 432258
rect 506942 432224 506976 432258
rect 507529 433114 507563 433148
rect 507619 433114 507653 433148
rect 507709 433114 507743 433148
rect 507799 433114 507833 433148
rect 507889 433114 507923 433148
rect 507979 433114 508013 433148
rect 508069 433114 508103 433148
rect 508159 433114 508193 433148
rect 508249 433114 508283 433148
rect 507416 433036 507450 433070
rect 507416 432946 507450 432980
rect 507416 432856 507450 432890
rect 507416 432766 507450 432800
rect 507416 432676 507450 432710
rect 507416 432586 507450 432620
rect 507416 432496 507450 432530
rect 507416 432406 507450 432440
rect 507416 432316 507450 432350
rect 508306 433002 508340 433036
rect 508306 432912 508340 432946
rect 508306 432822 508340 432856
rect 508306 432732 508340 432766
rect 508306 432642 508340 432676
rect 508306 432552 508340 432586
rect 508306 432462 508340 432496
rect 508306 432372 508340 432406
rect 508306 432282 508340 432316
rect 507510 432224 507544 432258
rect 507600 432224 507634 432258
rect 507690 432224 507724 432258
rect 507780 432224 507814 432258
rect 507870 432224 507904 432258
rect 507960 432224 507994 432258
rect 508050 432224 508084 432258
rect 508140 432224 508174 432258
rect 508230 432224 508264 432258
rect 508817 433114 508851 433148
rect 508907 433114 508941 433148
rect 508997 433114 509031 433148
rect 509087 433114 509121 433148
rect 509177 433114 509211 433148
rect 509267 433114 509301 433148
rect 509357 433114 509391 433148
rect 509447 433114 509481 433148
rect 509537 433114 509571 433148
rect 508704 433036 508738 433070
rect 508704 432946 508738 432980
rect 508704 432856 508738 432890
rect 508704 432766 508738 432800
rect 508704 432676 508738 432710
rect 508704 432586 508738 432620
rect 508704 432496 508738 432530
rect 508704 432406 508738 432440
rect 508704 432316 508738 432350
rect 509594 433002 509628 433036
rect 509594 432912 509628 432946
rect 509594 432822 509628 432856
rect 509594 432732 509628 432766
rect 509594 432642 509628 432676
rect 509594 432552 509628 432586
rect 509594 432462 509628 432496
rect 509594 432372 509628 432406
rect 509594 432282 509628 432316
rect 508798 432224 508832 432258
rect 508888 432224 508922 432258
rect 508978 432224 509012 432258
rect 509068 432224 509102 432258
rect 509158 432224 509192 432258
rect 509248 432224 509282 432258
rect 509338 432224 509372 432258
rect 509428 432224 509462 432258
rect 509518 432224 509552 432258
rect 510105 433114 510139 433148
rect 510195 433114 510229 433148
rect 510285 433114 510319 433148
rect 510375 433114 510409 433148
rect 510465 433114 510499 433148
rect 510555 433114 510589 433148
rect 510645 433114 510679 433148
rect 510735 433114 510769 433148
rect 510825 433114 510859 433148
rect 509992 433036 510026 433070
rect 509992 432946 510026 432980
rect 509992 432856 510026 432890
rect 509992 432766 510026 432800
rect 509992 432676 510026 432710
rect 509992 432586 510026 432620
rect 509992 432496 510026 432530
rect 509992 432406 510026 432440
rect 509992 432316 510026 432350
rect 510882 433002 510916 433036
rect 510882 432912 510916 432946
rect 510882 432822 510916 432856
rect 510882 432732 510916 432766
rect 510882 432642 510916 432676
rect 510882 432552 510916 432586
rect 510882 432462 510916 432496
rect 510882 432372 510916 432406
rect 510882 432282 510916 432316
rect 510086 432224 510120 432258
rect 510176 432224 510210 432258
rect 510266 432224 510300 432258
rect 510356 432224 510390 432258
rect 510446 432224 510480 432258
rect 510536 432224 510570 432258
rect 510626 432224 510660 432258
rect 510716 432224 510750 432258
rect 510806 432224 510840 432258
rect 511393 433114 511427 433148
rect 511483 433114 511517 433148
rect 511573 433114 511607 433148
rect 511663 433114 511697 433148
rect 511753 433114 511787 433148
rect 511843 433114 511877 433148
rect 511933 433114 511967 433148
rect 512023 433114 512057 433148
rect 512113 433114 512147 433148
rect 511280 433036 511314 433070
rect 511280 432946 511314 432980
rect 511280 432856 511314 432890
rect 511280 432766 511314 432800
rect 511280 432676 511314 432710
rect 511280 432586 511314 432620
rect 511280 432496 511314 432530
rect 511280 432406 511314 432440
rect 511280 432316 511314 432350
rect 512170 433002 512204 433036
rect 512170 432912 512204 432946
rect 512170 432822 512204 432856
rect 512170 432732 512204 432766
rect 512170 432642 512204 432676
rect 512170 432552 512204 432586
rect 512170 432462 512204 432496
rect 512170 432372 512204 432406
rect 512170 432282 512204 432316
rect 511374 432224 511408 432258
rect 511464 432224 511498 432258
rect 511554 432224 511588 432258
rect 511644 432224 511678 432258
rect 511734 432224 511768 432258
rect 511824 432224 511858 432258
rect 511914 432224 511948 432258
rect 512004 432224 512038 432258
rect 512094 432224 512128 432258
rect 512681 433114 512715 433148
rect 512771 433114 512805 433148
rect 512861 433114 512895 433148
rect 512951 433114 512985 433148
rect 513041 433114 513075 433148
rect 513131 433114 513165 433148
rect 513221 433114 513255 433148
rect 513311 433114 513345 433148
rect 513401 433114 513435 433148
rect 512568 433036 512602 433070
rect 512568 432946 512602 432980
rect 512568 432856 512602 432890
rect 512568 432766 512602 432800
rect 512568 432676 512602 432710
rect 512568 432586 512602 432620
rect 512568 432496 512602 432530
rect 512568 432406 512602 432440
rect 512568 432316 512602 432350
rect 513458 433002 513492 433036
rect 513458 432912 513492 432946
rect 513458 432822 513492 432856
rect 513458 432732 513492 432766
rect 513458 432642 513492 432676
rect 513458 432552 513492 432586
rect 513458 432462 513492 432496
rect 513458 432372 513492 432406
rect 513458 432282 513492 432316
rect 512662 432224 512696 432258
rect 512752 432224 512786 432258
rect 512842 432224 512876 432258
rect 512932 432224 512966 432258
rect 513022 432224 513056 432258
rect 513112 432224 513146 432258
rect 513202 432224 513236 432258
rect 513292 432224 513326 432258
rect 513382 432224 513416 432258
rect 562252 455178 567482 455212
rect 562156 454013 562190 455115
rect 567544 454013 567578 455115
rect 562252 453916 567482 453950
<< poly >>
rect 562316 495402 562516 495428
rect 562574 495402 562774 495428
rect 562832 495402 563032 495428
rect 563090 495402 563290 495428
rect 563348 495402 563548 495428
rect 563606 495402 563806 495428
rect 563864 495402 564064 495428
rect 564122 495402 564322 495428
rect 564380 495402 564580 495428
rect 564638 495402 564838 495428
rect 564896 495402 565096 495428
rect 565154 495402 565354 495428
rect 565412 495402 565612 495428
rect 565670 495402 565870 495428
rect 565928 495402 566128 495428
rect 566186 495402 566386 495428
rect 566444 495402 566644 495428
rect 566702 495402 566902 495428
rect 566960 495402 567160 495428
rect 567218 495402 567418 495428
rect 562316 494355 562516 494402
rect 562316 494321 562332 494355
rect 562500 494321 562516 494355
rect 562316 494305 562516 494321
rect 562574 494355 562774 494402
rect 562574 494321 562590 494355
rect 562758 494321 562774 494355
rect 562574 494305 562774 494321
rect 562832 494355 563032 494402
rect 562832 494321 562848 494355
rect 563016 494321 563032 494355
rect 562832 494305 563032 494321
rect 563090 494355 563290 494402
rect 563090 494321 563106 494355
rect 563274 494321 563290 494355
rect 563090 494305 563290 494321
rect 563348 494355 563548 494402
rect 563348 494321 563364 494355
rect 563532 494321 563548 494355
rect 563348 494305 563548 494321
rect 563606 494355 563806 494402
rect 563606 494321 563622 494355
rect 563790 494321 563806 494355
rect 563606 494305 563806 494321
rect 563864 494355 564064 494402
rect 563864 494321 563880 494355
rect 564048 494321 564064 494355
rect 563864 494305 564064 494321
rect 564122 494355 564322 494402
rect 564122 494321 564138 494355
rect 564306 494321 564322 494355
rect 564122 494305 564322 494321
rect 564380 494355 564580 494402
rect 564380 494321 564396 494355
rect 564564 494321 564580 494355
rect 564380 494305 564580 494321
rect 564638 494355 564838 494402
rect 564638 494321 564654 494355
rect 564822 494321 564838 494355
rect 564638 494305 564838 494321
rect 564896 494355 565096 494402
rect 564896 494321 564912 494355
rect 565080 494321 565096 494355
rect 564896 494305 565096 494321
rect 565154 494355 565354 494402
rect 565154 494321 565170 494355
rect 565338 494321 565354 494355
rect 565154 494305 565354 494321
rect 565412 494355 565612 494402
rect 565412 494321 565428 494355
rect 565596 494321 565612 494355
rect 565412 494305 565612 494321
rect 565670 494355 565870 494402
rect 565670 494321 565686 494355
rect 565854 494321 565870 494355
rect 565670 494305 565870 494321
rect 565928 494355 566128 494402
rect 565928 494321 565944 494355
rect 566112 494321 566128 494355
rect 565928 494305 566128 494321
rect 566186 494355 566386 494402
rect 566186 494321 566202 494355
rect 566370 494321 566386 494355
rect 566186 494305 566386 494321
rect 566444 494355 566644 494402
rect 566444 494321 566460 494355
rect 566628 494321 566644 494355
rect 566444 494305 566644 494321
rect 566702 494355 566902 494402
rect 566702 494321 566718 494355
rect 566886 494321 566902 494355
rect 566702 494305 566902 494321
rect 566960 494355 567160 494402
rect 566960 494321 566976 494355
rect 567144 494321 567160 494355
rect 566960 494305 567160 494321
rect 567218 494355 567418 494402
rect 567218 494321 567234 494355
rect 567402 494321 567418 494355
rect 567218 494305 567418 494321
rect 572476 495436 572676 495462
rect 572734 495436 572934 495462
rect 572992 495436 573192 495462
rect 573250 495436 573450 495462
rect 573508 495436 573708 495462
rect 573766 495436 573966 495462
rect 574024 495436 574224 495462
rect 574282 495436 574482 495462
rect 574540 495436 574740 495462
rect 574798 495436 574998 495462
rect 575056 495436 575256 495462
rect 575314 495436 575514 495462
rect 575572 495436 575772 495462
rect 575830 495436 576030 495462
rect 576088 495436 576288 495462
rect 576346 495436 576546 495462
rect 576604 495436 576804 495462
rect 576862 495436 577062 495462
rect 577120 495436 577320 495462
rect 577378 495436 577578 495462
rect 572476 494398 572676 494436
rect 572476 494364 572492 494398
rect 572660 494364 572676 494398
rect 572476 494348 572676 494364
rect 572734 494398 572934 494436
rect 572734 494364 572750 494398
rect 572918 494364 572934 494398
rect 572734 494348 572934 494364
rect 572992 494398 573192 494436
rect 572992 494364 573008 494398
rect 573176 494364 573192 494398
rect 572992 494348 573192 494364
rect 573250 494398 573450 494436
rect 573250 494364 573266 494398
rect 573434 494364 573450 494398
rect 573250 494348 573450 494364
rect 573508 494398 573708 494436
rect 573508 494364 573524 494398
rect 573692 494364 573708 494398
rect 573508 494348 573708 494364
rect 573766 494398 573966 494436
rect 573766 494364 573782 494398
rect 573950 494364 573966 494398
rect 573766 494348 573966 494364
rect 574024 494398 574224 494436
rect 574024 494364 574040 494398
rect 574208 494364 574224 494398
rect 574024 494348 574224 494364
rect 574282 494398 574482 494436
rect 574282 494364 574298 494398
rect 574466 494364 574482 494398
rect 574282 494348 574482 494364
rect 574540 494398 574740 494436
rect 574540 494364 574556 494398
rect 574724 494364 574740 494398
rect 574540 494348 574740 494364
rect 574798 494398 574998 494436
rect 574798 494364 574814 494398
rect 574982 494364 574998 494398
rect 574798 494348 574998 494364
rect 575056 494398 575256 494436
rect 575056 494364 575072 494398
rect 575240 494364 575256 494398
rect 575056 494348 575256 494364
rect 575314 494398 575514 494436
rect 575314 494364 575330 494398
rect 575498 494364 575514 494398
rect 575314 494348 575514 494364
rect 575572 494398 575772 494436
rect 575572 494364 575588 494398
rect 575756 494364 575772 494398
rect 575572 494348 575772 494364
rect 575830 494398 576030 494436
rect 575830 494364 575846 494398
rect 576014 494364 576030 494398
rect 575830 494348 576030 494364
rect 576088 494398 576288 494436
rect 576088 494364 576104 494398
rect 576272 494364 576288 494398
rect 576088 494348 576288 494364
rect 576346 494398 576546 494436
rect 576346 494364 576362 494398
rect 576530 494364 576546 494398
rect 576346 494348 576546 494364
rect 576604 494398 576804 494436
rect 576604 494364 576620 494398
rect 576788 494364 576804 494398
rect 576604 494348 576804 494364
rect 576862 494398 577062 494436
rect 576862 494364 576878 494398
rect 577046 494364 577062 494398
rect 576862 494348 577062 494364
rect 577120 494398 577320 494436
rect 577120 494364 577136 494398
rect 577304 494364 577320 494398
rect 577120 494348 577320 494364
rect 577378 494398 577578 494436
rect 577378 494364 577394 494398
rect 577562 494364 577578 494398
rect 577378 494348 577578 494364
rect 506532 472318 506558 472718
rect 506958 472702 507046 472718
rect 506958 472334 506996 472702
rect 507030 472334 507046 472702
rect 506958 472318 507046 472334
rect 506532 471860 506558 472260
rect 506958 472244 507046 472260
rect 506958 471876 506996 472244
rect 507030 471876 507046 472244
rect 506958 471860 507046 471876
rect 506532 471402 506558 471802
rect 506958 471786 507046 471802
rect 506958 471418 506996 471786
rect 507030 471418 507046 471786
rect 506958 471402 507046 471418
rect 506532 470944 506558 471344
rect 506958 471328 507046 471344
rect 506958 470960 506996 471328
rect 507030 470960 507046 471328
rect 506958 470944 507046 470960
rect 506532 470486 506558 470886
rect 506958 470870 507046 470886
rect 506958 470502 506996 470870
rect 507030 470502 507046 470870
rect 506958 470486 507046 470502
rect 506532 470028 506558 470428
rect 506958 470412 507046 470428
rect 506958 470044 506996 470412
rect 507030 470044 507046 470412
rect 506958 470028 507046 470044
rect 503062 469114 503088 469514
rect 505668 469498 505765 469514
rect 505668 469130 505715 469498
rect 505749 469130 505765 469498
rect 505668 469114 505765 469130
rect 503062 468542 503088 468942
rect 505668 468926 505765 468942
rect 505668 468558 505715 468926
rect 505749 468558 505765 468926
rect 505668 468542 505765 468558
rect 503062 467970 503088 468370
rect 505668 468354 505765 468370
rect 505668 467986 505715 468354
rect 505749 467986 505765 468354
rect 509832 468200 510232 468216
rect 509832 468166 509848 468200
rect 510216 468166 510232 468200
rect 509832 468128 510232 468166
rect 505668 467970 505765 467986
rect 503062 467398 503088 467798
rect 505668 467782 505765 467798
rect 505668 467414 505715 467782
rect 505749 467414 505765 467782
rect 505668 467398 505765 467414
rect 506254 467388 506280 467788
rect 508080 467772 508168 467788
rect 508080 467404 508118 467772
rect 508152 467404 508168 467772
rect 508080 467388 508168 467404
rect 503062 466826 503088 467226
rect 505668 467210 505765 467226
rect 505668 466842 505715 467210
rect 505749 466842 505765 467210
rect 505668 466826 505765 466842
rect 506254 466816 506280 467216
rect 508080 467200 508168 467216
rect 508080 466832 508118 467200
rect 508152 466832 508168 467200
rect 508080 466816 508168 466832
rect 503062 466254 503088 466654
rect 505668 466638 505765 466654
rect 505668 466270 505715 466638
rect 505749 466270 505765 466638
rect 505668 466254 505765 466270
rect 506254 466244 506280 466644
rect 508080 466628 508168 466644
rect 508080 466260 508118 466628
rect 508152 466260 508168 466628
rect 508080 466244 508168 466260
rect 503062 465682 503088 466082
rect 505668 466066 505765 466082
rect 505668 465698 505715 466066
rect 505749 465698 505765 466066
rect 505668 465682 505765 465698
rect 506254 465672 506280 466072
rect 508080 466056 508168 466072
rect 508080 465688 508118 466056
rect 508152 465688 508168 466056
rect 508080 465672 508168 465688
rect 503062 465110 503088 465510
rect 505668 465494 505765 465510
rect 505668 465126 505715 465494
rect 505749 465126 505765 465494
rect 505668 465110 505765 465126
rect 506254 465100 506280 465500
rect 508080 465484 508168 465500
rect 508080 465116 508118 465484
rect 508152 465116 508168 465484
rect 508080 465100 508168 465116
rect 503062 464538 503088 464938
rect 505668 464922 505765 464938
rect 505668 464554 505715 464922
rect 505749 464554 505765 464922
rect 505668 464538 505765 464554
rect 506254 464528 506280 464928
rect 508080 464912 508168 464928
rect 508080 464544 508118 464912
rect 508152 464544 508168 464912
rect 508080 464528 508168 464544
rect 503062 463966 503088 464366
rect 505668 464350 505765 464366
rect 505668 463982 505715 464350
rect 505749 463982 505765 464350
rect 505668 463966 505765 463982
rect 506254 463956 506280 464356
rect 508080 464340 508168 464356
rect 508080 463972 508118 464340
rect 508152 463972 508168 464340
rect 508080 463956 508168 463972
rect 503062 463394 503088 463794
rect 505668 463778 505765 463794
rect 505668 463410 505715 463778
rect 505749 463410 505765 463778
rect 505668 463394 505765 463410
rect 506254 463384 506280 463784
rect 508080 463768 508168 463784
rect 508080 463400 508118 463768
rect 508152 463400 508168 463768
rect 508080 463384 508168 463400
rect 503062 462822 503088 463222
rect 505668 463206 505765 463222
rect 505668 462838 505715 463206
rect 505749 462838 505765 463206
rect 505668 462822 505765 462838
rect 509832 462702 510232 462728
rect 503062 462250 503088 462650
rect 505668 462634 505765 462650
rect 505668 462266 505715 462634
rect 505749 462266 505765 462634
rect 505668 462250 505765 462266
rect 503062 461678 503088 462078
rect 505668 462062 505765 462078
rect 505668 461694 505715 462062
rect 505749 461694 505765 462062
rect 505668 461678 505765 461694
rect 503029 459690 503126 459706
rect 503029 459322 503045 459690
rect 503079 459322 503126 459690
rect 503029 459306 503126 459322
rect 510866 459306 510892 459706
rect 503029 459232 503126 459248
rect 503029 458864 503045 459232
rect 503079 458864 503126 459232
rect 503029 458848 503126 458864
rect 510866 458848 510892 459248
rect 503029 458774 503126 458790
rect 503029 458406 503045 458774
rect 503079 458406 503126 458774
rect 503029 458390 503126 458406
rect 510866 458390 510892 458790
rect 503029 458316 503126 458332
rect 503029 457948 503045 458316
rect 503079 457948 503126 458316
rect 503029 457932 503126 457948
rect 510866 457932 510892 458332
rect 503029 457858 503126 457874
rect 503029 457490 503045 457858
rect 503079 457490 503126 457858
rect 503029 457474 503126 457490
rect 510866 457474 510892 457874
rect 503029 457400 503126 457416
rect 503029 457032 503045 457400
rect 503079 457032 503126 457400
rect 503029 457016 503126 457032
rect 510866 457016 510892 457416
rect 503029 456942 503126 456958
rect 503029 456574 503045 456942
rect 503079 456574 503126 456942
rect 503029 456558 503126 456574
rect 510866 456558 510892 456958
rect 503029 456484 503126 456500
rect 503029 456116 503045 456484
rect 503079 456116 503126 456484
rect 503029 456100 503126 456116
rect 510866 456100 510892 456500
rect 503029 456026 503126 456042
rect 503029 455658 503045 456026
rect 503079 455658 503126 456026
rect 503029 455642 503126 455658
rect 510866 455642 510892 456042
rect 503029 455568 503126 455584
rect 503029 455200 503045 455568
rect 503079 455200 503126 455568
rect 503029 455184 503126 455200
rect 510866 455184 510892 455584
rect 503029 455110 503126 455126
rect 503029 454742 503045 455110
rect 503079 454742 503126 455110
rect 503029 454726 503126 454742
rect 510866 454726 510892 455126
rect 503029 453732 503126 453748
rect 503029 453364 503045 453732
rect 503079 453364 503126 453732
rect 503029 453348 503126 453364
rect 510866 453348 510892 453748
rect 503029 453274 503126 453290
rect 503029 452906 503045 453274
rect 503079 452906 503126 453274
rect 503029 452890 503126 452906
rect 510866 452890 510892 453290
rect 503029 452816 503126 452832
rect 503029 452448 503045 452816
rect 503079 452448 503126 452816
rect 503029 452432 503126 452448
rect 510866 452432 510892 452832
rect 503029 452358 503126 452374
rect 503029 451990 503045 452358
rect 503079 451990 503126 452358
rect 503029 451974 503126 451990
rect 510866 451974 510892 452374
rect 503029 451900 503126 451916
rect 503029 451532 503045 451900
rect 503079 451532 503126 451900
rect 503029 451516 503126 451532
rect 510866 451516 510892 451916
rect 503029 451442 503126 451458
rect 503029 451074 503045 451442
rect 503079 451074 503126 451442
rect 503029 451058 503126 451074
rect 510866 451058 510892 451458
rect 503029 450984 503126 451000
rect 503029 450616 503045 450984
rect 503079 450616 503126 450984
rect 503029 450600 503126 450616
rect 510866 450600 510892 451000
rect 503029 450526 503126 450542
rect 503029 450158 503045 450526
rect 503079 450158 503126 450526
rect 503029 450142 503126 450158
rect 510866 450142 510892 450542
rect 503029 450068 503126 450084
rect 503029 449700 503045 450068
rect 503079 449700 503126 450068
rect 503029 449684 503126 449700
rect 510866 449684 510892 450084
rect 503029 449610 503126 449626
rect 503029 449242 503045 449610
rect 503079 449242 503126 449610
rect 503029 449226 503126 449242
rect 510866 449226 510892 449626
rect 503029 448232 503126 448248
rect 503029 447864 503045 448232
rect 503079 447864 503126 448232
rect 503029 447848 503126 447864
rect 510866 447848 510892 448248
rect 503029 447774 503126 447790
rect 503029 447406 503045 447774
rect 503079 447406 503126 447774
rect 503029 447390 503126 447406
rect 510866 447390 510892 447790
rect 503029 447316 503126 447332
rect 503029 446948 503045 447316
rect 503079 446948 503126 447316
rect 503029 446932 503126 446948
rect 510866 446932 510892 447332
rect 503029 446858 503126 446874
rect 503029 446490 503045 446858
rect 503079 446490 503126 446858
rect 503029 446474 503126 446490
rect 510866 446474 510892 446874
rect 503029 446400 503126 446416
rect 503029 446032 503045 446400
rect 503079 446032 503126 446400
rect 503029 446016 503126 446032
rect 510866 446016 510892 446416
rect 503029 445942 503126 445958
rect 503029 445574 503045 445942
rect 503079 445574 503126 445942
rect 503029 445558 503126 445574
rect 510866 445558 510892 445958
rect 503029 445484 503126 445500
rect 503029 445116 503045 445484
rect 503079 445116 503126 445484
rect 503029 445100 503126 445116
rect 510866 445100 510892 445500
rect 503029 445026 503126 445042
rect 503029 444658 503045 445026
rect 503079 444658 503126 445026
rect 503029 444642 503126 444658
rect 510866 444642 510892 445042
rect 503029 444568 503126 444584
rect 503029 444200 503045 444568
rect 503079 444200 503126 444568
rect 503029 444184 503126 444200
rect 510866 444184 510892 444584
rect 503029 444110 503126 444126
rect 503029 443742 503045 444110
rect 503079 443742 503126 444110
rect 503029 443726 503126 443742
rect 510866 443726 510892 444126
rect 503029 443652 503126 443668
rect 503029 443284 503045 443652
rect 503079 443284 503126 443652
rect 503029 443268 503126 443284
rect 510866 443268 510892 443668
rect 562316 455100 562516 455126
rect 562574 455100 562774 455126
rect 562832 455100 563032 455126
rect 563090 455100 563290 455126
rect 563348 455100 563548 455126
rect 563606 455100 563806 455126
rect 563864 455100 564064 455126
rect 564122 455100 564322 455126
rect 564380 455100 564580 455126
rect 564638 455100 564838 455126
rect 564896 455100 565096 455126
rect 565154 455100 565354 455126
rect 565412 455100 565612 455126
rect 565670 455100 565870 455126
rect 565928 455100 566128 455126
rect 566186 455100 566386 455126
rect 566444 455100 566644 455126
rect 566702 455100 566902 455126
rect 566960 455100 567160 455126
rect 567218 455100 567418 455126
rect 562316 454053 562516 454100
rect 562316 454019 562332 454053
rect 562500 454019 562516 454053
rect 562316 454003 562516 454019
rect 562574 454053 562774 454100
rect 562574 454019 562590 454053
rect 562758 454019 562774 454053
rect 562574 454003 562774 454019
rect 562832 454053 563032 454100
rect 562832 454019 562848 454053
rect 563016 454019 563032 454053
rect 562832 454003 563032 454019
rect 563090 454053 563290 454100
rect 563090 454019 563106 454053
rect 563274 454019 563290 454053
rect 563090 454003 563290 454019
rect 563348 454053 563548 454100
rect 563348 454019 563364 454053
rect 563532 454019 563548 454053
rect 563348 454003 563548 454019
rect 563606 454053 563806 454100
rect 563606 454019 563622 454053
rect 563790 454019 563806 454053
rect 563606 454003 563806 454019
rect 563864 454053 564064 454100
rect 563864 454019 563880 454053
rect 564048 454019 564064 454053
rect 563864 454003 564064 454019
rect 564122 454053 564322 454100
rect 564122 454019 564138 454053
rect 564306 454019 564322 454053
rect 564122 454003 564322 454019
rect 564380 454053 564580 454100
rect 564380 454019 564396 454053
rect 564564 454019 564580 454053
rect 564380 454003 564580 454019
rect 564638 454053 564838 454100
rect 564638 454019 564654 454053
rect 564822 454019 564838 454053
rect 564638 454003 564838 454019
rect 564896 454053 565096 454100
rect 564896 454019 564912 454053
rect 565080 454019 565096 454053
rect 564896 454003 565096 454019
rect 565154 454053 565354 454100
rect 565154 454019 565170 454053
rect 565338 454019 565354 454053
rect 565154 454003 565354 454019
rect 565412 454053 565612 454100
rect 565412 454019 565428 454053
rect 565596 454019 565612 454053
rect 565412 454003 565612 454019
rect 565670 454053 565870 454100
rect 565670 454019 565686 454053
rect 565854 454019 565870 454053
rect 565670 454003 565870 454019
rect 565928 454053 566128 454100
rect 565928 454019 565944 454053
rect 566112 454019 566128 454053
rect 565928 454003 566128 454019
rect 566186 454053 566386 454100
rect 566186 454019 566202 454053
rect 566370 454019 566386 454053
rect 566186 454003 566386 454019
rect 566444 454053 566644 454100
rect 566444 454019 566460 454053
rect 566628 454019 566644 454053
rect 566444 454003 566644 454019
rect 566702 454053 566902 454100
rect 566702 454019 566718 454053
rect 566886 454019 566902 454053
rect 566702 454003 566902 454019
rect 566960 454053 567160 454100
rect 566960 454019 566976 454053
rect 567144 454019 567160 454053
rect 566960 454003 567160 454019
rect 567218 454053 567418 454100
rect 567218 454019 567234 454053
rect 567402 454019 567418 454053
rect 567218 454003 567418 454019
rect 572476 455134 572676 455160
rect 572734 455134 572934 455160
rect 572992 455134 573192 455160
rect 573250 455134 573450 455160
rect 573508 455134 573708 455160
rect 573766 455134 573966 455160
rect 574024 455134 574224 455160
rect 574282 455134 574482 455160
rect 574540 455134 574740 455160
rect 574798 455134 574998 455160
rect 575056 455134 575256 455160
rect 575314 455134 575514 455160
rect 575572 455134 575772 455160
rect 575830 455134 576030 455160
rect 576088 455134 576288 455160
rect 576346 455134 576546 455160
rect 576604 455134 576804 455160
rect 576862 455134 577062 455160
rect 577120 455134 577320 455160
rect 577378 455134 577578 455160
rect 572476 454096 572676 454134
rect 572476 454062 572492 454096
rect 572660 454062 572676 454096
rect 572476 454046 572676 454062
rect 572734 454096 572934 454134
rect 572734 454062 572750 454096
rect 572918 454062 572934 454096
rect 572734 454046 572934 454062
rect 572992 454096 573192 454134
rect 572992 454062 573008 454096
rect 573176 454062 573192 454096
rect 572992 454046 573192 454062
rect 573250 454096 573450 454134
rect 573250 454062 573266 454096
rect 573434 454062 573450 454096
rect 573250 454046 573450 454062
rect 573508 454096 573708 454134
rect 573508 454062 573524 454096
rect 573692 454062 573708 454096
rect 573508 454046 573708 454062
rect 573766 454096 573966 454134
rect 573766 454062 573782 454096
rect 573950 454062 573966 454096
rect 573766 454046 573966 454062
rect 574024 454096 574224 454134
rect 574024 454062 574040 454096
rect 574208 454062 574224 454096
rect 574024 454046 574224 454062
rect 574282 454096 574482 454134
rect 574282 454062 574298 454096
rect 574466 454062 574482 454096
rect 574282 454046 574482 454062
rect 574540 454096 574740 454134
rect 574540 454062 574556 454096
rect 574724 454062 574740 454096
rect 574540 454046 574740 454062
rect 574798 454096 574998 454134
rect 574798 454062 574814 454096
rect 574982 454062 574998 454096
rect 574798 454046 574998 454062
rect 575056 454096 575256 454134
rect 575056 454062 575072 454096
rect 575240 454062 575256 454096
rect 575056 454046 575256 454062
rect 575314 454096 575514 454134
rect 575314 454062 575330 454096
rect 575498 454062 575514 454096
rect 575314 454046 575514 454062
rect 575572 454096 575772 454134
rect 575572 454062 575588 454096
rect 575756 454062 575772 454096
rect 575572 454046 575772 454062
rect 575830 454096 576030 454134
rect 575830 454062 575846 454096
rect 576014 454062 576030 454096
rect 575830 454046 576030 454062
rect 576088 454096 576288 454134
rect 576088 454062 576104 454096
rect 576272 454062 576288 454096
rect 576088 454046 576288 454062
rect 576346 454096 576546 454134
rect 576346 454062 576362 454096
rect 576530 454062 576546 454096
rect 576346 454046 576546 454062
rect 576604 454096 576804 454134
rect 576604 454062 576620 454096
rect 576788 454062 576804 454096
rect 576604 454046 576804 454062
rect 576862 454096 577062 454134
rect 576862 454062 576878 454096
rect 577046 454062 577062 454096
rect 576862 454046 577062 454062
rect 577120 454096 577320 454134
rect 577120 454062 577136 454096
rect 577304 454062 577320 454096
rect 577120 454046 577320 454062
rect 577378 454096 577578 454134
rect 577378 454062 577394 454096
rect 577562 454062 577578 454096
rect 577378 454046 577578 454062
<< polycont >>
rect 562332 494321 562500 494355
rect 562590 494321 562758 494355
rect 562848 494321 563016 494355
rect 563106 494321 563274 494355
rect 563364 494321 563532 494355
rect 563622 494321 563790 494355
rect 563880 494321 564048 494355
rect 564138 494321 564306 494355
rect 564396 494321 564564 494355
rect 564654 494321 564822 494355
rect 564912 494321 565080 494355
rect 565170 494321 565338 494355
rect 565428 494321 565596 494355
rect 565686 494321 565854 494355
rect 565944 494321 566112 494355
rect 566202 494321 566370 494355
rect 566460 494321 566628 494355
rect 566718 494321 566886 494355
rect 566976 494321 567144 494355
rect 567234 494321 567402 494355
rect 572492 494364 572660 494398
rect 572750 494364 572918 494398
rect 573008 494364 573176 494398
rect 573266 494364 573434 494398
rect 573524 494364 573692 494398
rect 573782 494364 573950 494398
rect 574040 494364 574208 494398
rect 574298 494364 574466 494398
rect 574556 494364 574724 494398
rect 574814 494364 574982 494398
rect 575072 494364 575240 494398
rect 575330 494364 575498 494398
rect 575588 494364 575756 494398
rect 575846 494364 576014 494398
rect 576104 494364 576272 494398
rect 576362 494364 576530 494398
rect 576620 494364 576788 494398
rect 576878 494364 577046 494398
rect 577136 494364 577304 494398
rect 577394 494364 577562 494398
rect 506996 472334 507030 472702
rect 506996 471876 507030 472244
rect 506996 471418 507030 471786
rect 506996 470960 507030 471328
rect 506996 470502 507030 470870
rect 506996 470044 507030 470412
rect 505715 469130 505749 469498
rect 505715 468558 505749 468926
rect 505715 467986 505749 468354
rect 509848 468166 510216 468200
rect 505715 467414 505749 467782
rect 508118 467404 508152 467772
rect 505715 466842 505749 467210
rect 508118 466832 508152 467200
rect 505715 466270 505749 466638
rect 508118 466260 508152 466628
rect 505715 465698 505749 466066
rect 508118 465688 508152 466056
rect 505715 465126 505749 465494
rect 508118 465116 508152 465484
rect 505715 464554 505749 464922
rect 508118 464544 508152 464912
rect 505715 463982 505749 464350
rect 508118 463972 508152 464340
rect 505715 463410 505749 463778
rect 508118 463400 508152 463768
rect 505715 462838 505749 463206
rect 505715 462266 505749 462634
rect 505715 461694 505749 462062
rect 503045 459322 503079 459690
rect 503045 458864 503079 459232
rect 503045 458406 503079 458774
rect 503045 457948 503079 458316
rect 503045 457490 503079 457858
rect 503045 457032 503079 457400
rect 503045 456574 503079 456942
rect 503045 456116 503079 456484
rect 503045 455658 503079 456026
rect 503045 455200 503079 455568
rect 503045 454742 503079 455110
rect 503045 453364 503079 453732
rect 503045 452906 503079 453274
rect 503045 452448 503079 452816
rect 503045 451990 503079 452358
rect 503045 451532 503079 451900
rect 503045 451074 503079 451442
rect 503045 450616 503079 450984
rect 503045 450158 503079 450526
rect 503045 449700 503079 450068
rect 503045 449242 503079 449610
rect 503045 447864 503079 448232
rect 503045 447406 503079 447774
rect 503045 446948 503079 447316
rect 503045 446490 503079 446858
rect 503045 446032 503079 446400
rect 503045 445574 503079 445942
rect 503045 445116 503079 445484
rect 503045 444658 503079 445026
rect 503045 444200 503079 444568
rect 503045 443742 503079 444110
rect 503045 443284 503079 443652
rect 562332 454019 562500 454053
rect 562590 454019 562758 454053
rect 562848 454019 563016 454053
rect 563106 454019 563274 454053
rect 563364 454019 563532 454053
rect 563622 454019 563790 454053
rect 563880 454019 564048 454053
rect 564138 454019 564306 454053
rect 564396 454019 564564 454053
rect 564654 454019 564822 454053
rect 564912 454019 565080 454053
rect 565170 454019 565338 454053
rect 565428 454019 565596 454053
rect 565686 454019 565854 454053
rect 565944 454019 566112 454053
rect 566202 454019 566370 454053
rect 566460 454019 566628 454053
rect 566718 454019 566886 454053
rect 566976 454019 567144 454053
rect 567234 454019 567402 454053
rect 572492 454062 572660 454096
rect 572750 454062 572918 454096
rect 573008 454062 573176 454096
rect 573266 454062 573434 454096
rect 573524 454062 573692 454096
rect 573782 454062 573950 454096
rect 574040 454062 574208 454096
rect 574298 454062 574466 454096
rect 574556 454062 574724 454096
rect 574814 454062 574982 454096
rect 575072 454062 575240 454096
rect 575330 454062 575498 454096
rect 575588 454062 575756 454096
rect 575846 454062 576014 454096
rect 576104 454062 576272 454096
rect 576362 454062 576530 454096
rect 576620 454062 576788 454096
rect 576878 454062 577046 454096
rect 577136 454062 577304 454096
rect 577394 454062 577562 454096
<< xpolycontact >>
rect 517846 459314 518278 459884
rect 521602 459314 522034 459884
rect 517846 458496 518278 459066
rect 521602 458496 522034 459066
rect 517846 457678 518278 458248
rect 521602 457678 522034 458248
rect 518256 456042 518688 456612
rect 522988 456042 523420 456612
rect 518256 455224 518688 455794
rect 522988 455224 523420 455794
rect 518256 454406 518688 454976
rect 522988 454406 523420 454976
rect 518256 453588 518688 454158
rect 522988 453588 523420 454158
rect 516190 451134 516622 451704
rect 522926 451134 523358 451704
rect 516190 450316 516622 450886
rect 522926 450316 523358 450886
rect 516190 449498 516622 450068
rect 522926 449498 523358 450068
rect 516190 448680 516622 449250
rect 522926 448680 523358 449250
rect 516190 447862 516622 448432
rect 522926 447862 523358 448432
rect 516190 447044 516622 447614
rect 522926 447044 523358 447614
rect 516190 446226 516622 446796
rect 522926 446226 523358 446796
rect 516190 445408 516622 445978
rect 522926 445408 523358 445978
rect 516190 444590 516622 445160
rect 522926 444590 523358 445160
rect 516190 443772 516622 444342
rect 522926 443772 523358 444342
rect 516190 442954 516622 443524
rect 522926 442954 523358 443524
rect 516190 442136 516622 442706
rect 522926 442136 523358 442706
rect 516190 441318 516622 441888
rect 522926 441318 523358 441888
rect 516190 440500 516622 441070
rect 522926 440500 523358 441070
rect 516190 439682 516622 440252
rect 522926 439682 523358 440252
rect 516190 438864 516622 439434
rect 522926 438864 523358 439434
rect 516190 438046 516622 438616
rect 522926 438046 523358 438616
<< xpolyres >>
rect 518278 459314 521602 459884
rect 518278 458496 521602 459066
rect 518278 457678 521602 458248
rect 518688 456042 522988 456612
rect 518688 455224 522988 455794
rect 518688 454406 522988 454976
rect 518688 453588 522988 454158
rect 516622 451134 522926 451704
rect 516622 450316 522926 450886
rect 516622 449498 522926 450068
rect 516622 448680 522926 449250
rect 516622 447862 522926 448432
rect 516622 447044 522926 447614
rect 516622 446226 522926 446796
rect 516622 445408 522926 445978
rect 516622 444590 522926 445160
rect 516622 443772 522926 444342
rect 516622 442954 522926 443524
rect 516622 442136 522926 442706
rect 516622 441318 522926 441888
rect 516622 440500 522926 441070
rect 516622 439682 522926 440252
rect 516622 438864 522926 439434
rect 516622 438046 522926 438616
<< locali >>
rect 562156 495417 562190 495514
rect 567544 495417 567578 495514
rect 562270 495390 562304 495406
rect 562270 494398 562304 494414
rect 562528 495390 562562 495406
rect 562528 494355 562562 494414
rect 562786 495390 562820 495406
rect 562786 494398 562820 494414
rect 563044 495390 563078 495406
rect 563044 494355 563078 494414
rect 563302 495390 563336 495406
rect 563302 494398 563336 494414
rect 563560 495390 563594 495406
rect 563560 494355 563594 494414
rect 563818 495390 563852 495406
rect 563818 494398 563852 494414
rect 564076 495390 564110 495406
rect 564076 494355 564110 494414
rect 564334 495390 564368 495406
rect 564334 494398 564368 494414
rect 564592 495390 564626 495406
rect 564592 494355 564626 494414
rect 564850 495390 564884 495406
rect 564850 494398 564884 494414
rect 565108 495390 565142 495406
rect 565108 494355 565142 494414
rect 565366 495390 565400 495406
rect 565366 494398 565400 494414
rect 565624 495390 565658 495406
rect 565624 494355 565658 494414
rect 565882 495390 565916 495406
rect 565882 494398 565916 494414
rect 566140 495390 566174 495406
rect 566140 494355 566174 494414
rect 566398 495390 566432 495406
rect 566398 494398 566432 494414
rect 566656 495390 566690 495406
rect 566656 494355 566690 494414
rect 566914 495390 566948 495406
rect 566914 494398 566948 494414
rect 567172 495390 567206 495406
rect 567172 494355 567206 494414
rect 567430 495390 567464 495406
rect 567430 494398 567464 494414
rect 562270 494321 562332 494355
rect 562500 494321 562590 494355
rect 562758 494321 562848 494355
rect 563016 494321 563106 494355
rect 563274 494321 563364 494355
rect 563532 494321 563622 494355
rect 563790 494321 563880 494355
rect 564048 494321 564138 494355
rect 564306 494321 564396 494355
rect 564564 494321 564654 494355
rect 564822 494321 564912 494355
rect 565080 494321 565170 494355
rect 565338 494321 565428 494355
rect 565596 494321 565686 494355
rect 565854 494321 565944 494355
rect 566112 494321 566202 494355
rect 566370 494321 566460 494355
rect 566628 494321 566718 494355
rect 566886 494321 566976 494355
rect 567144 494321 567234 494355
rect 567402 494321 567464 494355
rect 562156 494252 562190 494315
rect 567544 494252 567578 494315
rect 572316 495452 572350 495548
rect 577704 495452 577738 495548
rect 572430 495424 572464 495440
rect 572430 494432 572464 494448
rect 572688 495424 572722 495440
rect 572688 494398 572722 494448
rect 572946 495424 572980 495440
rect 572946 494432 572980 494448
rect 573204 495424 573238 495440
rect 573204 494398 573238 494448
rect 573462 495424 573496 495440
rect 573462 494432 573496 494448
rect 573720 495424 573754 495440
rect 573720 494398 573754 494448
rect 573978 495424 574012 495440
rect 573978 494432 574012 494448
rect 574236 495424 574270 495440
rect 574236 494398 574270 494448
rect 574494 495424 574528 495440
rect 574494 494432 574528 494448
rect 574752 495424 574786 495440
rect 574752 494398 574786 494448
rect 575010 495424 575044 495440
rect 575010 494432 575044 494448
rect 575268 495424 575302 495440
rect 575268 494398 575302 494448
rect 575526 495424 575560 495440
rect 575526 494432 575560 494448
rect 575784 495424 575818 495440
rect 575784 494398 575818 494448
rect 576042 495424 576076 495440
rect 576042 494432 576076 494448
rect 576300 495424 576334 495440
rect 576300 494398 576334 494448
rect 576558 495424 576592 495440
rect 576558 494432 576592 494448
rect 576816 495424 576850 495440
rect 576816 494398 576850 494448
rect 577074 495424 577108 495440
rect 577074 494432 577108 494448
rect 577332 495424 577366 495440
rect 577332 494398 577366 494448
rect 577590 495424 577624 495440
rect 577590 494432 577624 494448
rect 572429 494364 572492 494398
rect 572660 494364 572750 494398
rect 572918 494364 573008 494398
rect 573176 494364 573266 494398
rect 573434 494364 573524 494398
rect 573692 494364 573782 494398
rect 573950 494364 574040 494398
rect 574208 494364 574298 494398
rect 574466 494364 574556 494398
rect 574724 494364 574814 494398
rect 574982 494364 575072 494398
rect 575240 494364 575330 494398
rect 575498 494364 575588 494398
rect 575756 494364 575846 494398
rect 576014 494364 576104 494398
rect 576272 494364 576362 494398
rect 576530 494364 576620 494398
rect 576788 494364 576878 494398
rect 577046 494364 577136 494398
rect 577304 494364 577394 494398
rect 577562 494364 577626 494398
rect 572316 494296 572350 494358
rect 577704 494296 577738 494358
rect 572316 494262 572412 494296
rect 577642 494262 577738 494296
rect 562156 494218 562252 494252
rect 567482 494218 567578 494252
rect 500320 475332 528616 475356
rect 500320 475308 527592 475332
rect 500320 474332 500368 475308
rect 500352 433044 500368 474332
rect 501368 475306 527592 475308
rect 501368 475284 503920 475306
rect 504020 475284 504144 475306
rect 504244 475284 504368 475306
rect 504468 475284 504592 475306
rect 504692 475284 504816 475306
rect 504916 475284 505040 475306
rect 505140 475284 505264 475306
rect 505364 475284 505488 475306
rect 505588 475284 505712 475306
rect 505812 475284 505936 475306
rect 506036 475284 506160 475306
rect 506260 475284 506384 475306
rect 506484 475284 506608 475306
rect 506708 475284 506832 475306
rect 506932 475284 507056 475306
rect 507156 475284 507280 475306
rect 507380 475284 507504 475306
rect 507604 475284 507728 475306
rect 507828 475284 507952 475306
rect 508052 475284 508176 475306
rect 508276 475284 508400 475306
rect 508500 475284 508624 475306
rect 508724 475284 508848 475306
rect 508948 475284 509072 475306
rect 509172 475284 509296 475306
rect 509396 475284 509520 475306
rect 509620 475284 509744 475306
rect 509844 475284 509968 475306
rect 510068 475284 510192 475306
rect 510292 475284 510416 475306
rect 510516 475284 517320 475306
rect 517420 475284 517544 475306
rect 517644 475284 517768 475306
rect 517868 475284 517992 475306
rect 518092 475284 518216 475306
rect 518316 475284 518440 475306
rect 518540 475284 518664 475306
rect 518764 475284 518888 475306
rect 518988 475284 519112 475306
rect 519212 475284 519336 475306
rect 519436 475284 519560 475306
rect 519660 475284 519784 475306
rect 519884 475284 520008 475306
rect 520108 475284 520232 475306
rect 520332 475284 520456 475306
rect 520556 475284 520680 475306
rect 520780 475284 520904 475306
rect 521004 475284 521128 475306
rect 521228 475284 521352 475306
rect 521452 475284 521576 475306
rect 521676 475284 521800 475306
rect 521900 475284 522024 475306
rect 522124 475284 522248 475306
rect 522348 475284 522472 475306
rect 522572 475284 522696 475306
rect 522796 475284 522920 475306
rect 523020 475284 523144 475306
rect 523244 475284 523368 475306
rect 523468 475284 523592 475306
rect 523692 475284 523816 475306
rect 523916 475284 527592 475306
rect 501368 474332 502392 475284
rect 501368 474280 501384 474332
rect 502376 474284 502392 474332
rect 526544 474332 527592 475284
rect 526544 474284 526560 474332
rect 502376 474268 526560 474284
rect 501368 474056 501384 474180
rect 501368 473832 501384 473956
rect 501368 473608 501384 473732
rect 501368 473384 501384 473508
rect 501368 473160 501384 473284
rect 506516 473256 507124 473272
rect 501368 472936 501384 473060
rect 506516 472856 506532 473256
rect 507108 472856 507124 473256
rect 506516 472840 507124 472856
rect 501368 472712 501384 472836
rect 506554 472764 507030 472840
rect 506554 472730 506570 472764
rect 506946 472730 507030 472764
rect 506996 472702 507030 472730
rect 501368 472488 501384 472612
rect 501368 472264 501384 472388
rect 506996 472318 507030 472334
rect 506554 472272 506570 472306
rect 506946 472272 506962 472306
rect 506996 472244 507030 472260
rect 501368 472040 501384 472164
rect 501368 471816 501384 471940
rect 506554 471814 506570 471848
rect 506946 471814 506962 471848
rect 506996 471786 507030 471876
rect 501368 471592 501384 471716
rect 501368 471368 501384 471492
rect 506554 471356 506570 471390
rect 506946 471356 506962 471390
rect 506996 471328 507030 471418
rect 501368 471144 501384 471268
rect 501368 470920 501384 471044
rect 506554 470898 506570 470932
rect 506946 470898 506962 470932
rect 506996 470870 507030 470960
rect 501368 470696 501384 470820
rect 507082 471870 507278 471886
rect 507082 471858 507186 471870
rect 507082 471806 507094 471858
rect 507146 471806 507186 471858
rect 507082 470942 507186 471806
rect 507082 470890 507094 470942
rect 507146 470890 507186 470942
rect 507082 470878 507186 470890
rect 507262 470878 507278 471870
rect 507082 470862 507278 470878
rect 501368 470472 501384 470596
rect 506996 470486 507030 470502
rect 506554 470440 506570 470474
rect 506946 470440 506962 470474
rect 506996 470412 507030 470428
rect 501368 470248 501384 470372
rect 503210 470202 505580 470218
rect 501368 470024 501384 470148
rect 503210 470102 503226 470202
rect 505568 470102 505580 470202
rect 503210 470086 505580 470102
rect 506996 470016 507030 470044
rect 506554 469982 506570 470016
rect 506946 469982 507030 470016
rect 501368 469800 501384 469924
rect 506554 469906 507030 469982
rect 506516 469890 507124 469906
rect 501368 469576 501384 469700
rect 503084 469526 503100 469560
rect 505656 469526 505672 469560
rect 505715 469498 505749 469514
rect 501368 469352 501384 469476
rect 506516 469490 506532 469890
rect 507108 469490 507124 469890
rect 506516 469474 507124 469490
rect 501368 469128 501384 469252
rect 505715 469114 505749 469130
rect 503084 469068 503100 469102
rect 505656 469068 505672 469102
rect 501368 468904 501384 469028
rect 503084 468954 503100 468988
rect 505656 468954 505672 468988
rect 505715 468926 505749 468942
rect 501368 468680 501384 468804
rect 501368 468456 501384 468580
rect 505715 468542 505749 468558
rect 510460 468840 510824 468850
rect 503084 468496 503100 468530
rect 505656 468496 505672 468530
rect 503084 468382 503100 468416
rect 505656 468382 505672 468416
rect 506452 468386 508084 468402
rect 501368 468232 501384 468356
rect 505715 468354 505749 468370
rect 506452 468286 506468 468386
rect 508068 468286 508084 468386
rect 506452 468270 508084 468286
rect 501368 468008 501384 468132
rect 509832 468166 509848 468200
rect 510216 468166 510232 468200
rect 505715 467970 505749 467986
rect 509786 468116 509820 468132
rect 503084 467924 503100 467958
rect 505656 467924 505672 467958
rect 501368 467784 501384 467908
rect 503084 467810 503100 467844
rect 505656 467810 505672 467844
rect 506276 467800 506292 467834
rect 508068 467800 508084 467834
rect 505715 467782 505749 467798
rect 501368 463810 501384 467684
rect 505715 467398 505749 467414
rect 508118 467772 508152 467788
rect 508118 467388 508152 467404
rect 503084 467352 503100 467386
rect 505656 467352 505672 467386
rect 506276 467342 506292 467376
rect 508068 467342 508084 467376
rect 503084 467238 503100 467272
rect 505656 467238 505672 467272
rect 506276 467228 506292 467262
rect 508068 467228 508084 467262
rect 505715 467210 505749 467226
rect 505715 466826 505749 466842
rect 508118 467200 508152 467216
rect 508118 466816 508152 466832
rect 503084 466780 503100 466814
rect 505656 466780 505672 466814
rect 506276 466770 506292 466804
rect 508068 466770 508084 466804
rect 503084 466666 503100 466700
rect 505656 466666 505672 466700
rect 506276 466656 506292 466690
rect 508068 466656 508084 466690
rect 505715 466638 505749 466654
rect 502606 466620 502738 466632
rect 502606 464278 502622 466620
rect 502722 464278 502738 466620
rect 505715 466254 505749 466270
rect 508118 466628 508152 466644
rect 508118 466244 508152 466260
rect 503084 466208 503100 466242
rect 505656 466208 505672 466242
rect 506276 466198 506292 466232
rect 508068 466198 508084 466232
rect 503084 466094 503100 466128
rect 505656 466094 505672 466128
rect 506276 466084 506292 466118
rect 508068 466084 508084 466118
rect 505715 466066 505749 466082
rect 505715 465682 505749 465698
rect 508118 466056 508152 466072
rect 508118 465672 508152 465688
rect 503084 465636 503100 465670
rect 505656 465636 505672 465670
rect 506276 465626 506292 465660
rect 508068 465626 508084 465660
rect 503084 465522 503100 465556
rect 505656 465522 505672 465556
rect 506276 465512 506292 465546
rect 508068 465512 508084 465546
rect 505715 465494 505749 465510
rect 505715 465110 505749 465126
rect 508118 465484 508152 465500
rect 508118 465100 508152 465116
rect 503084 465064 503100 465098
rect 505656 465064 505672 465098
rect 506276 465054 506292 465088
rect 508068 465054 508084 465088
rect 503084 464950 503100 464984
rect 505656 464950 505672 464984
rect 506276 464940 506292 464974
rect 508068 464940 508084 464974
rect 505715 464922 505749 464938
rect 505715 464538 505749 464554
rect 508118 464912 508152 464928
rect 508118 464528 508152 464544
rect 503084 464492 503100 464526
rect 505656 464492 505672 464526
rect 506276 464482 506292 464516
rect 508068 464482 508084 464516
rect 503084 464378 503100 464412
rect 505656 464378 505672 464412
rect 506276 464368 506292 464402
rect 508068 464368 508084 464402
rect 502606 464262 502738 464278
rect 505715 464350 505749 464366
rect 505715 463966 505749 463982
rect 508118 464340 508152 464356
rect 508118 463956 508152 463972
rect 503084 463920 503100 463954
rect 505656 463920 505672 463954
rect 506276 463910 506292 463944
rect 508068 463910 508084 463944
rect 503084 463806 503100 463840
rect 505656 463806 505672 463840
rect 506276 463796 506292 463830
rect 508068 463796 508084 463830
rect 505715 463778 505749 463794
rect 501368 463586 501384 463710
rect 501368 463362 501384 463486
rect 505715 463394 505749 463410
rect 508118 463768 508152 463784
rect 508118 463384 508152 463400
rect 503084 463348 503100 463382
rect 505656 463348 505672 463382
rect 506276 463338 506292 463372
rect 508068 463338 508084 463372
rect 501368 463138 501384 463262
rect 503084 463234 503100 463268
rect 505656 463234 505672 463268
rect 505715 463206 505749 463222
rect 501368 462914 501384 463038
rect 505715 462822 505749 462838
rect 506452 462886 508084 462902
rect 501368 462690 501384 462814
rect 503084 462776 503100 462810
rect 505656 462776 505672 462810
rect 506452 462786 506468 462886
rect 508068 462786 508084 462886
rect 506452 462770 508084 462786
rect 509786 462724 509820 462740
rect 510244 468116 510278 468132
rect 510244 462724 510278 462740
rect 503084 462662 503100 462696
rect 505656 462662 505672 462696
rect 505715 462634 505749 462650
rect 501368 462466 501384 462590
rect 501368 462242 501384 462366
rect 510460 462376 510470 468840
rect 510814 462376 510824 468840
rect 510460 462366 510824 462376
rect 505715 462250 505749 462266
rect 503084 462204 503100 462238
rect 505656 462204 505672 462238
rect 501368 462018 501384 462142
rect 503084 462090 503100 462124
rect 505656 462090 505672 462124
rect 505715 462062 505749 462078
rect 501368 461794 501384 461918
rect 501368 461570 501384 461694
rect 505715 461678 505749 461694
rect 503084 461632 503100 461666
rect 505656 461632 505672 461666
rect 501368 461346 501384 461470
rect 501368 461122 501384 461246
rect 503210 461074 505580 461090
rect 501368 460898 501384 461022
rect 503210 460974 503226 461074
rect 505568 460974 505580 461074
rect 503210 460958 505580 460974
rect 501368 460674 501384 460798
rect 517028 460724 517532 460728
rect 521592 460724 522034 460734
rect 516606 460708 522942 460724
rect 501368 460450 501384 460574
rect 502428 460352 510728 460452
rect 501368 460226 501384 460350
rect 501368 460002 501384 460126
rect 502428 459952 502528 460352
rect 502628 460252 510728 460352
rect 502628 460052 503528 460252
rect 510528 460052 510728 460252
rect 516606 460138 516622 460708
rect 522926 460138 522942 460708
rect 516606 460122 522942 460138
rect 502628 459952 510728 460052
rect 501368 459778 501384 459902
rect 502428 459852 510728 459952
rect 517028 459884 517532 460122
rect 521592 459884 522034 460122
rect 503122 459718 503138 459752
rect 510854 459718 510870 459752
rect 503045 459690 503079 459706
rect 501368 459554 501384 459678
rect 501368 459330 501384 459454
rect 503045 459306 503079 459322
rect 517028 459314 517846 459884
rect 521592 459314 521602 459884
rect 503122 459260 503138 459294
rect 510854 459260 510870 459294
rect 503045 459232 503079 459248
rect 501368 459106 501384 459230
rect 501368 458882 501384 459006
rect 503045 458848 503079 458864
rect 503122 458802 503138 458836
rect 510854 458802 510870 458836
rect 501368 458658 501384 458782
rect 503045 458774 503079 458790
rect 501368 458434 501384 458558
rect 503045 458390 503079 458406
rect 503122 458344 503138 458378
rect 510854 458344 510870 458378
rect 501368 458210 501384 458334
rect 503045 458316 503079 458332
rect 501368 457986 501384 458110
rect 503045 457932 503079 457948
rect 503122 457886 503138 457920
rect 510854 457886 510870 457920
rect 501368 457762 501384 457886
rect 503045 457858 503079 457874
rect 501368 457538 501384 457662
rect 503045 457474 503079 457490
rect 517028 457480 517536 459314
rect 521592 459066 522034 459314
rect 521592 458496 521602 459066
rect 521592 458248 522034 458496
rect 517846 457480 518278 457678
rect 521592 457678 521602 458248
rect 521592 457480 522034 457678
rect 522430 457480 523420 457486
rect 516606 457464 523420 457480
rect 501368 457314 501384 457438
rect 503122 457428 503138 457462
rect 510854 457428 510870 457462
rect 503045 457400 503079 457416
rect 501368 437540 501384 457214
rect 503045 457016 503079 457032
rect 503122 456970 503138 457004
rect 510854 456970 510870 457004
rect 503045 456942 503079 456958
rect 516606 456894 516622 457464
rect 522926 456894 523420 457464
rect 516606 456882 523420 456894
rect 516606 456878 522942 456882
rect 517028 456868 517536 456878
rect 503045 456558 503079 456574
rect 518158 456612 518684 456878
rect 522988 456612 523420 456882
rect 503122 456512 503138 456546
rect 510854 456512 510870 456546
rect 503045 456484 503079 456500
rect 503045 456100 503079 456116
rect 503122 456054 503138 456088
rect 510854 456054 510870 456088
rect 518158 456042 518256 456612
rect 503045 456026 503079 456042
rect 518158 455936 518688 456042
rect 503045 455642 503079 455658
rect 503122 455596 503138 455630
rect 510854 455596 510870 455630
rect 503045 455568 503079 455584
rect 503045 455184 503079 455200
rect 503122 455138 503138 455172
rect 510854 455138 510870 455172
rect 503045 455110 503079 455126
rect 503045 454726 503079 454742
rect 503122 454680 503138 454714
rect 510854 454680 510870 454714
rect 502428 454442 510728 454542
rect 502428 454042 502528 454442
rect 502628 454342 510728 454442
rect 502628 454142 503528 454342
rect 510528 454142 510728 454342
rect 502628 454042 510728 454142
rect 502428 453942 510728 454042
rect 518158 454158 518688 454274
rect 503122 453760 503138 453794
rect 510854 453760 510870 453794
rect 503045 453732 503079 453748
rect 503045 453348 503079 453364
rect 518158 453588 518256 454158
rect 503122 453302 503138 453336
rect 510854 453302 510870 453336
rect 503045 453274 503079 453290
rect 503045 452890 503079 452906
rect 503122 452844 503138 452878
rect 510854 452844 510870 452878
rect 503045 452816 503079 452832
rect 503045 452432 503079 452448
rect 516190 452520 516622 452528
rect 518158 452520 518688 453588
rect 522926 453588 522988 454158
rect 522926 452520 523420 453588
rect 516190 452504 523420 452520
rect 503122 452386 503138 452420
rect 510854 452386 510870 452420
rect 503045 452358 503079 452374
rect 503045 451974 503079 451990
rect 503122 451928 503138 451962
rect 510854 451928 510870 451962
rect 516190 451934 516622 452504
rect 522926 451934 523420 452504
rect 516190 451918 523420 451934
rect 503045 451900 503079 451916
rect 503045 451516 503079 451532
rect 516190 451704 516622 451918
rect 503122 451470 503138 451504
rect 510854 451470 510870 451504
rect 503045 451442 503079 451458
rect 522926 451704 523420 451918
rect 523358 451134 523420 451704
rect 503045 451058 503079 451074
rect 503122 451012 503138 451046
rect 510854 451012 510870 451046
rect 503045 450984 503079 451000
rect 503045 450600 503079 450616
rect 503122 450554 503138 450588
rect 510854 450554 510870 450588
rect 503045 450526 503079 450542
rect 503045 450142 503079 450158
rect 503122 450096 503138 450130
rect 510854 450096 510870 450130
rect 503045 450068 503079 450084
rect 503045 449684 503079 449700
rect 503122 449638 503138 449672
rect 510854 449638 510870 449672
rect 503045 449610 503079 449626
rect 503045 449226 503079 449242
rect 503122 449180 503138 449214
rect 510854 449180 510870 449214
rect 502428 448942 510728 449042
rect 502428 448542 502528 448942
rect 502628 448842 510728 448942
rect 502628 448642 503528 448842
rect 510528 448642 510728 448842
rect 502628 448542 510728 448642
rect 502428 448442 510728 448542
rect 503122 448260 503138 448294
rect 510854 448260 510870 448294
rect 503045 448232 503079 448248
rect 503045 447848 503079 447864
rect 503122 447802 503138 447836
rect 510854 447802 510870 447836
rect 503045 447774 503079 447790
rect 503045 447390 503079 447406
rect 503122 447344 503138 447378
rect 510854 447344 510870 447378
rect 503045 447316 503079 447332
rect 503045 446932 503079 446948
rect 503122 446886 503138 446920
rect 510854 446886 510870 446920
rect 503045 446858 503079 446874
rect 503045 446474 503079 446490
rect 503122 446428 503138 446462
rect 510854 446428 510870 446462
rect 503045 446400 503079 446416
rect 503045 446016 503079 446032
rect 503122 445970 503138 446004
rect 510854 445970 510870 446004
rect 503045 445942 503079 445958
rect 503045 445558 503079 445574
rect 503122 445512 503138 445546
rect 510854 445512 510870 445546
rect 503045 445484 503079 445500
rect 503045 445100 503079 445116
rect 503122 445054 503138 445088
rect 510854 445054 510870 445088
rect 503045 445026 503079 445042
rect 503045 444642 503079 444658
rect 503122 444596 503138 444630
rect 510854 444596 510870 444630
rect 503045 444568 503079 444584
rect 503045 444184 503079 444200
rect 503122 444138 503138 444172
rect 510854 444138 510870 444172
rect 503045 444110 503079 444126
rect 503045 443726 503079 443742
rect 503122 443680 503138 443714
rect 510854 443680 510870 443714
rect 503045 443652 503079 443668
rect 503045 443268 503079 443284
rect 503122 443222 503138 443256
rect 510854 443222 510870 443256
rect 502426 442986 510726 443086
rect 502426 442586 502526 442986
rect 502626 442886 510726 442986
rect 502626 442686 503526 442886
rect 510526 442686 510726 442886
rect 502626 442586 510726 442686
rect 502426 442486 510726 442586
rect 503370 438448 513674 438482
rect 503370 438414 503486 438448
rect 503520 438414 503576 438448
rect 503610 438414 503666 438448
rect 503700 438414 503756 438448
rect 503790 438414 503846 438448
rect 503880 438414 503936 438448
rect 503970 438414 504026 438448
rect 504060 438414 504116 438448
rect 504150 438414 504206 438448
rect 504240 438414 504296 438448
rect 504330 438414 504386 438448
rect 504420 438414 504476 438448
rect 504510 438414 504566 438448
rect 504600 438414 504774 438448
rect 504808 438414 504864 438448
rect 504898 438414 504954 438448
rect 504988 438414 505044 438448
rect 505078 438414 505134 438448
rect 505168 438414 505224 438448
rect 505258 438414 505314 438448
rect 505348 438414 505404 438448
rect 505438 438414 505494 438448
rect 505528 438414 505584 438448
rect 505618 438414 505674 438448
rect 505708 438414 505764 438448
rect 505798 438414 505854 438448
rect 505888 438414 506062 438448
rect 506096 438414 506152 438448
rect 506186 438414 506242 438448
rect 506276 438414 506332 438448
rect 506366 438414 506422 438448
rect 506456 438414 506512 438448
rect 506546 438414 506602 438448
rect 506636 438414 506692 438448
rect 506726 438414 506782 438448
rect 506816 438414 506872 438448
rect 506906 438414 506962 438448
rect 506996 438414 507052 438448
rect 507086 438414 507142 438448
rect 507176 438414 507350 438448
rect 507384 438414 507440 438448
rect 507474 438414 507530 438448
rect 507564 438414 507620 438448
rect 507654 438414 507710 438448
rect 507744 438414 507800 438448
rect 507834 438414 507890 438448
rect 507924 438414 507980 438448
rect 508014 438414 508070 438448
rect 508104 438414 508160 438448
rect 508194 438414 508250 438448
rect 508284 438414 508340 438448
rect 508374 438414 508430 438448
rect 508464 438414 508638 438448
rect 508672 438414 508728 438448
rect 508762 438414 508818 438448
rect 508852 438414 508908 438448
rect 508942 438414 508998 438448
rect 509032 438414 509088 438448
rect 509122 438414 509178 438448
rect 509212 438414 509268 438448
rect 509302 438414 509358 438448
rect 509392 438414 509448 438448
rect 509482 438414 509538 438448
rect 509572 438414 509628 438448
rect 509662 438414 509718 438448
rect 509752 438414 509926 438448
rect 509960 438414 510016 438448
rect 510050 438414 510106 438448
rect 510140 438414 510196 438448
rect 510230 438414 510286 438448
rect 510320 438414 510376 438448
rect 510410 438414 510466 438448
rect 510500 438414 510556 438448
rect 510590 438414 510646 438448
rect 510680 438414 510736 438448
rect 510770 438414 510826 438448
rect 510860 438414 510916 438448
rect 510950 438414 511006 438448
rect 511040 438414 511214 438448
rect 511248 438414 511304 438448
rect 511338 438414 511394 438448
rect 511428 438414 511484 438448
rect 511518 438414 511574 438448
rect 511608 438414 511664 438448
rect 511698 438414 511754 438448
rect 511788 438414 511844 438448
rect 511878 438414 511934 438448
rect 511968 438414 512024 438448
rect 512058 438414 512114 438448
rect 512148 438414 512204 438448
rect 512238 438414 512294 438448
rect 512328 438414 512502 438448
rect 512536 438414 512592 438448
rect 512626 438414 512682 438448
rect 512716 438414 512772 438448
rect 512806 438414 512862 438448
rect 512896 438414 512952 438448
rect 512986 438414 513042 438448
rect 513076 438414 513132 438448
rect 513166 438414 513222 438448
rect 513256 438414 513312 438448
rect 513346 438414 513402 438448
rect 513436 438414 513492 438448
rect 513526 438414 513582 438448
rect 513616 438414 513674 438448
rect 503370 438352 513674 438414
rect 503370 438318 503402 438352
rect 503436 438318 504589 438352
rect 504623 438318 504690 438352
rect 504724 438318 505877 438352
rect 505911 438318 505978 438352
rect 506012 438318 507165 438352
rect 507199 438318 507266 438352
rect 507300 438318 508453 438352
rect 508487 438318 508554 438352
rect 508588 438318 509741 438352
rect 509775 438318 509842 438352
rect 509876 438318 511029 438352
rect 511063 438318 511130 438352
rect 511164 438318 512317 438352
rect 512351 438318 512418 438352
rect 512452 438318 513605 438352
rect 513639 438318 513674 438352
rect 503370 438300 513674 438318
rect 503370 438266 503665 438300
rect 503699 438266 503755 438300
rect 503789 438266 503845 438300
rect 503879 438266 503935 438300
rect 503969 438266 504025 438300
rect 504059 438266 504115 438300
rect 504149 438266 504205 438300
rect 504239 438266 504295 438300
rect 504329 438266 504385 438300
rect 504419 438266 504953 438300
rect 504987 438266 505043 438300
rect 505077 438266 505133 438300
rect 505167 438266 505223 438300
rect 505257 438266 505313 438300
rect 505347 438266 505403 438300
rect 505437 438266 505493 438300
rect 505527 438266 505583 438300
rect 505617 438266 505673 438300
rect 505707 438266 506241 438300
rect 506275 438266 506331 438300
rect 506365 438266 506421 438300
rect 506455 438266 506511 438300
rect 506545 438266 506601 438300
rect 506635 438266 506691 438300
rect 506725 438266 506781 438300
rect 506815 438266 506871 438300
rect 506905 438266 506961 438300
rect 506995 438266 507529 438300
rect 507563 438266 507619 438300
rect 507653 438266 507709 438300
rect 507743 438266 507799 438300
rect 507833 438266 507889 438300
rect 507923 438266 507979 438300
rect 508013 438266 508069 438300
rect 508103 438266 508159 438300
rect 508193 438266 508249 438300
rect 508283 438266 508817 438300
rect 508851 438266 508907 438300
rect 508941 438266 508997 438300
rect 509031 438266 509087 438300
rect 509121 438266 509177 438300
rect 509211 438266 509267 438300
rect 509301 438266 509357 438300
rect 509391 438266 509447 438300
rect 509481 438266 509537 438300
rect 509571 438266 510105 438300
rect 510139 438266 510195 438300
rect 510229 438266 510285 438300
rect 510319 438266 510375 438300
rect 510409 438266 510465 438300
rect 510499 438266 510555 438300
rect 510589 438266 510645 438300
rect 510679 438266 510735 438300
rect 510769 438266 510825 438300
rect 510859 438266 511393 438300
rect 511427 438266 511483 438300
rect 511517 438266 511573 438300
rect 511607 438266 511663 438300
rect 511697 438266 511753 438300
rect 511787 438266 511843 438300
rect 511877 438266 511933 438300
rect 511967 438266 512023 438300
rect 512057 438266 512113 438300
rect 512147 438266 512681 438300
rect 512715 438266 512771 438300
rect 512805 438266 512861 438300
rect 512895 438266 512951 438300
rect 512985 438266 513041 438300
rect 513075 438266 513131 438300
rect 513165 438266 513221 438300
rect 513255 438266 513311 438300
rect 513345 438266 513401 438300
rect 513435 438266 513674 438300
rect 503370 438262 513674 438266
rect 503370 438228 503402 438262
rect 503436 438247 504589 438262
rect 503436 438228 503605 438247
rect 503370 438222 503605 438228
rect 503370 438188 503552 438222
rect 503586 438188 503605 438222
rect 503370 438172 503605 438188
rect 504423 438228 504589 438247
rect 504623 438228 504690 438262
rect 504724 438247 505877 438262
rect 504724 438228 504893 438247
rect 504423 438222 504893 438228
rect 504423 438188 504840 438222
rect 504874 438188 504893 438222
rect 503370 438138 503402 438172
rect 503436 438138 503605 438172
rect 503370 438132 503605 438138
rect 503370 438098 503552 438132
rect 503586 438098 503605 438132
rect 503370 438082 503605 438098
rect 503370 438048 503402 438082
rect 503436 438048 503605 438082
rect 503370 438042 503605 438048
rect 503370 438008 503552 438042
rect 503586 438008 503605 438042
rect 503370 437992 503605 438008
rect 503370 437958 503402 437992
rect 503436 437958 503605 437992
rect 503370 437952 503605 437958
rect 503370 437918 503552 437952
rect 503586 437918 503605 437952
rect 503370 437902 503605 437918
rect 503370 437868 503402 437902
rect 503436 437868 503605 437902
rect 503370 437862 503605 437868
rect 503370 437828 503552 437862
rect 503586 437828 503605 437862
rect 503370 437812 503605 437828
rect 503370 437778 503402 437812
rect 503436 437778 503605 437812
rect 503370 437772 503605 437778
rect 503370 437738 503552 437772
rect 503586 437738 503605 437772
rect 503370 437722 503605 437738
rect 503370 437688 503402 437722
rect 503436 437688 503605 437722
rect 503370 437682 503605 437688
rect 503370 437648 503552 437682
rect 503586 437648 503605 437682
rect 503370 437632 503605 437648
rect 503370 437598 503402 437632
rect 503436 437598 503605 437632
rect 503370 437592 503605 437598
rect 503370 437558 503552 437592
rect 503586 437558 503605 437592
rect 503370 437542 503605 437558
rect 503370 437508 503402 437542
rect 503436 437508 503605 437542
rect 503370 437502 503605 437508
rect 503370 437468 503552 437502
rect 503586 437468 503605 437502
rect 503667 438124 504361 438185
rect 503667 438090 503728 438124
rect 503762 438112 503818 438124
rect 503852 438112 503908 438124
rect 503942 438112 503998 438124
rect 503774 438090 503818 438112
rect 503874 438090 503908 438112
rect 503974 438090 503998 438112
rect 504032 438112 504088 438124
rect 504032 438090 504040 438112
rect 503667 438078 503740 438090
rect 503774 438078 503840 438090
rect 503874 438078 503940 438090
rect 503974 438078 504040 438090
rect 504074 438090 504088 438112
rect 504122 438112 504178 438124
rect 504122 438090 504140 438112
rect 504074 438078 504140 438090
rect 504174 438090 504178 438112
rect 504212 438112 504268 438124
rect 504212 438090 504240 438112
rect 504302 438090 504361 438124
rect 504174 438078 504240 438090
rect 504274 438078 504361 438090
rect 503667 438034 504361 438078
rect 503667 438000 503728 438034
rect 503762 438012 503818 438034
rect 503852 438012 503908 438034
rect 503942 438012 503998 438034
rect 503774 438000 503818 438012
rect 503874 438000 503908 438012
rect 503974 438000 503998 438012
rect 504032 438012 504088 438034
rect 504032 438000 504040 438012
rect 503667 437978 503740 438000
rect 503774 437978 503840 438000
rect 503874 437978 503940 438000
rect 503974 437978 504040 438000
rect 504074 438000 504088 438012
rect 504122 438012 504178 438034
rect 504122 438000 504140 438012
rect 504074 437978 504140 438000
rect 504174 438000 504178 438012
rect 504212 438012 504268 438034
rect 504212 438000 504240 438012
rect 504302 438000 504361 438034
rect 504174 437978 504240 438000
rect 504274 437978 504361 438000
rect 503667 437944 504361 437978
rect 503667 437910 503728 437944
rect 503762 437912 503818 437944
rect 503852 437912 503908 437944
rect 503942 437912 503998 437944
rect 503774 437910 503818 437912
rect 503874 437910 503908 437912
rect 503974 437910 503998 437912
rect 504032 437912 504088 437944
rect 504032 437910 504040 437912
rect 503667 437878 503740 437910
rect 503774 437878 503840 437910
rect 503874 437878 503940 437910
rect 503974 437878 504040 437910
rect 504074 437910 504088 437912
rect 504122 437912 504178 437944
rect 504122 437910 504140 437912
rect 504074 437878 504140 437910
rect 504174 437910 504178 437912
rect 504212 437912 504268 437944
rect 504212 437910 504240 437912
rect 504302 437910 504361 437944
rect 504174 437878 504240 437910
rect 504274 437878 504361 437910
rect 503667 437854 504361 437878
rect 503667 437820 503728 437854
rect 503762 437820 503818 437854
rect 503852 437820 503908 437854
rect 503942 437820 503998 437854
rect 504032 437820 504088 437854
rect 504122 437820 504178 437854
rect 504212 437820 504268 437854
rect 504302 437820 504361 437854
rect 503667 437812 504361 437820
rect 503667 437778 503740 437812
rect 503774 437778 503840 437812
rect 503874 437778 503940 437812
rect 503974 437778 504040 437812
rect 504074 437778 504140 437812
rect 504174 437778 504240 437812
rect 504274 437778 504361 437812
rect 503667 437764 504361 437778
rect 503667 437730 503728 437764
rect 503762 437730 503818 437764
rect 503852 437730 503908 437764
rect 503942 437730 503998 437764
rect 504032 437730 504088 437764
rect 504122 437730 504178 437764
rect 504212 437730 504268 437764
rect 504302 437730 504361 437764
rect 503667 437712 504361 437730
rect 503667 437678 503740 437712
rect 503774 437678 503840 437712
rect 503874 437678 503940 437712
rect 503974 437678 504040 437712
rect 504074 437678 504140 437712
rect 504174 437678 504240 437712
rect 504274 437678 504361 437712
rect 503667 437674 504361 437678
rect 503667 437640 503728 437674
rect 503762 437640 503818 437674
rect 503852 437640 503908 437674
rect 503942 437640 503998 437674
rect 504032 437640 504088 437674
rect 504122 437640 504178 437674
rect 504212 437640 504268 437674
rect 504302 437640 504361 437674
rect 503667 437612 504361 437640
rect 503667 437584 503740 437612
rect 503774 437584 503840 437612
rect 503874 437584 503940 437612
rect 503974 437584 504040 437612
rect 503667 437550 503728 437584
rect 503774 437578 503818 437584
rect 503874 437578 503908 437584
rect 503974 437578 503998 437584
rect 503762 437550 503818 437578
rect 503852 437550 503908 437578
rect 503942 437550 503998 437578
rect 504032 437578 504040 437584
rect 504074 437584 504140 437612
rect 504074 437578 504088 437584
rect 504032 437550 504088 437578
rect 504122 437578 504140 437584
rect 504174 437584 504240 437612
rect 504274 437584 504361 437612
rect 504174 437578 504178 437584
rect 504122 437550 504178 437578
rect 504212 437578 504240 437584
rect 504212 437550 504268 437578
rect 504302 437550 504361 437584
rect 503667 437491 504361 437550
rect 504423 438154 504442 438188
rect 504476 438172 504893 438188
rect 505711 438228 505877 438247
rect 505911 438228 505978 438262
rect 506012 438247 507165 438262
rect 506012 438228 506181 438247
rect 505711 438222 506181 438228
rect 505711 438188 506128 438222
rect 506162 438188 506181 438222
rect 504476 438154 504589 438172
rect 504423 438138 504589 438154
rect 504623 438138 504690 438172
rect 504724 438138 504893 438172
rect 504423 438132 504893 438138
rect 504423 438098 504840 438132
rect 504874 438098 504893 438132
rect 504423 438064 504442 438098
rect 504476 438082 504893 438098
rect 504476 438064 504589 438082
rect 504423 438048 504589 438064
rect 504623 438048 504690 438082
rect 504724 438048 504893 438082
rect 504423 438042 504893 438048
rect 504423 438008 504840 438042
rect 504874 438008 504893 438042
rect 504423 437974 504442 438008
rect 504476 437992 504893 438008
rect 504476 437974 504589 437992
rect 504423 437958 504589 437974
rect 504623 437958 504690 437992
rect 504724 437958 504893 437992
rect 504423 437952 504893 437958
rect 504423 437918 504840 437952
rect 504874 437918 504893 437952
rect 504423 437884 504442 437918
rect 504476 437902 504893 437918
rect 504476 437884 504589 437902
rect 504423 437868 504589 437884
rect 504623 437868 504690 437902
rect 504724 437868 504893 437902
rect 504423 437862 504893 437868
rect 504423 437828 504840 437862
rect 504874 437828 504893 437862
rect 504423 437794 504442 437828
rect 504476 437812 504893 437828
rect 504476 437794 504589 437812
rect 504423 437778 504589 437794
rect 504623 437778 504690 437812
rect 504724 437778 504893 437812
rect 504423 437772 504893 437778
rect 504423 437738 504840 437772
rect 504874 437738 504893 437772
rect 504423 437704 504442 437738
rect 504476 437722 504893 437738
rect 504476 437704 504589 437722
rect 504423 437688 504589 437704
rect 504623 437688 504690 437722
rect 504724 437688 504893 437722
rect 504423 437682 504893 437688
rect 504423 437648 504840 437682
rect 504874 437648 504893 437682
rect 504423 437614 504442 437648
rect 504476 437632 504893 437648
rect 504476 437614 504589 437632
rect 504423 437598 504589 437614
rect 504623 437598 504690 437632
rect 504724 437598 504893 437632
rect 504423 437592 504893 437598
rect 504423 437558 504840 437592
rect 504874 437558 504893 437592
rect 504423 437524 504442 437558
rect 504476 437542 504893 437558
rect 504476 437524 504589 437542
rect 504423 437508 504589 437524
rect 504623 437508 504690 437542
rect 504724 437508 504893 437542
rect 504423 437502 504893 437508
rect 503370 437452 503605 437468
rect 501368 437316 501384 437440
rect 503370 437418 503402 437452
rect 503436 437429 503605 437452
rect 504423 437468 504840 437502
rect 504874 437468 504893 437502
rect 504955 438124 505649 438185
rect 504955 438090 505016 438124
rect 505050 438112 505106 438124
rect 505140 438112 505196 438124
rect 505230 438112 505286 438124
rect 505062 438090 505106 438112
rect 505162 438090 505196 438112
rect 505262 438090 505286 438112
rect 505320 438112 505376 438124
rect 505320 438090 505328 438112
rect 504955 438078 505028 438090
rect 505062 438078 505128 438090
rect 505162 438078 505228 438090
rect 505262 438078 505328 438090
rect 505362 438090 505376 438112
rect 505410 438112 505466 438124
rect 505410 438090 505428 438112
rect 505362 438078 505428 438090
rect 505462 438090 505466 438112
rect 505500 438112 505556 438124
rect 505500 438090 505528 438112
rect 505590 438090 505649 438124
rect 505462 438078 505528 438090
rect 505562 438078 505649 438090
rect 504955 438034 505649 438078
rect 504955 438000 505016 438034
rect 505050 438012 505106 438034
rect 505140 438012 505196 438034
rect 505230 438012 505286 438034
rect 505062 438000 505106 438012
rect 505162 438000 505196 438012
rect 505262 438000 505286 438012
rect 505320 438012 505376 438034
rect 505320 438000 505328 438012
rect 504955 437978 505028 438000
rect 505062 437978 505128 438000
rect 505162 437978 505228 438000
rect 505262 437978 505328 438000
rect 505362 438000 505376 438012
rect 505410 438012 505466 438034
rect 505410 438000 505428 438012
rect 505362 437978 505428 438000
rect 505462 438000 505466 438012
rect 505500 438012 505556 438034
rect 505500 438000 505528 438012
rect 505590 438000 505649 438034
rect 505462 437978 505528 438000
rect 505562 437978 505649 438000
rect 504955 437944 505649 437978
rect 504955 437910 505016 437944
rect 505050 437912 505106 437944
rect 505140 437912 505196 437944
rect 505230 437912 505286 437944
rect 505062 437910 505106 437912
rect 505162 437910 505196 437912
rect 505262 437910 505286 437912
rect 505320 437912 505376 437944
rect 505320 437910 505328 437912
rect 504955 437878 505028 437910
rect 505062 437878 505128 437910
rect 505162 437878 505228 437910
rect 505262 437878 505328 437910
rect 505362 437910 505376 437912
rect 505410 437912 505466 437944
rect 505410 437910 505428 437912
rect 505362 437878 505428 437910
rect 505462 437910 505466 437912
rect 505500 437912 505556 437944
rect 505500 437910 505528 437912
rect 505590 437910 505649 437944
rect 505462 437878 505528 437910
rect 505562 437878 505649 437910
rect 504955 437854 505649 437878
rect 504955 437820 505016 437854
rect 505050 437820 505106 437854
rect 505140 437820 505196 437854
rect 505230 437820 505286 437854
rect 505320 437820 505376 437854
rect 505410 437820 505466 437854
rect 505500 437820 505556 437854
rect 505590 437820 505649 437854
rect 504955 437812 505649 437820
rect 504955 437778 505028 437812
rect 505062 437778 505128 437812
rect 505162 437778 505228 437812
rect 505262 437778 505328 437812
rect 505362 437778 505428 437812
rect 505462 437778 505528 437812
rect 505562 437778 505649 437812
rect 504955 437764 505649 437778
rect 504955 437730 505016 437764
rect 505050 437730 505106 437764
rect 505140 437730 505196 437764
rect 505230 437730 505286 437764
rect 505320 437730 505376 437764
rect 505410 437730 505466 437764
rect 505500 437730 505556 437764
rect 505590 437730 505649 437764
rect 504955 437712 505649 437730
rect 504955 437678 505028 437712
rect 505062 437678 505128 437712
rect 505162 437678 505228 437712
rect 505262 437678 505328 437712
rect 505362 437678 505428 437712
rect 505462 437678 505528 437712
rect 505562 437678 505649 437712
rect 504955 437674 505649 437678
rect 504955 437640 505016 437674
rect 505050 437640 505106 437674
rect 505140 437640 505196 437674
rect 505230 437640 505286 437674
rect 505320 437640 505376 437674
rect 505410 437640 505466 437674
rect 505500 437640 505556 437674
rect 505590 437640 505649 437674
rect 504955 437612 505649 437640
rect 504955 437584 505028 437612
rect 505062 437584 505128 437612
rect 505162 437584 505228 437612
rect 505262 437584 505328 437612
rect 504955 437550 505016 437584
rect 505062 437578 505106 437584
rect 505162 437578 505196 437584
rect 505262 437578 505286 437584
rect 505050 437550 505106 437578
rect 505140 437550 505196 437578
rect 505230 437550 505286 437578
rect 505320 437578 505328 437584
rect 505362 437584 505428 437612
rect 505362 437578 505376 437584
rect 505320 437550 505376 437578
rect 505410 437578 505428 437584
rect 505462 437584 505528 437612
rect 505562 437584 505649 437612
rect 505462 437578 505466 437584
rect 505410 437550 505466 437578
rect 505500 437578 505528 437584
rect 505500 437550 505556 437578
rect 505590 437550 505649 437584
rect 504955 437491 505649 437550
rect 505711 438154 505730 438188
rect 505764 438172 506181 438188
rect 506999 438228 507165 438247
rect 507199 438228 507266 438262
rect 507300 438247 508453 438262
rect 507300 438228 507469 438247
rect 506999 438222 507469 438228
rect 506999 438188 507416 438222
rect 507450 438188 507469 438222
rect 505764 438154 505877 438172
rect 505711 438138 505877 438154
rect 505911 438138 505978 438172
rect 506012 438138 506181 438172
rect 505711 438132 506181 438138
rect 505711 438098 506128 438132
rect 506162 438098 506181 438132
rect 505711 438064 505730 438098
rect 505764 438082 506181 438098
rect 505764 438064 505877 438082
rect 505711 438048 505877 438064
rect 505911 438048 505978 438082
rect 506012 438048 506181 438082
rect 505711 438042 506181 438048
rect 505711 438008 506128 438042
rect 506162 438008 506181 438042
rect 505711 437974 505730 438008
rect 505764 437992 506181 438008
rect 505764 437974 505877 437992
rect 505711 437958 505877 437974
rect 505911 437958 505978 437992
rect 506012 437958 506181 437992
rect 505711 437952 506181 437958
rect 505711 437918 506128 437952
rect 506162 437918 506181 437952
rect 505711 437884 505730 437918
rect 505764 437902 506181 437918
rect 505764 437884 505877 437902
rect 505711 437868 505877 437884
rect 505911 437868 505978 437902
rect 506012 437868 506181 437902
rect 505711 437862 506181 437868
rect 505711 437828 506128 437862
rect 506162 437828 506181 437862
rect 505711 437794 505730 437828
rect 505764 437812 506181 437828
rect 505764 437794 505877 437812
rect 505711 437778 505877 437794
rect 505911 437778 505978 437812
rect 506012 437778 506181 437812
rect 505711 437772 506181 437778
rect 505711 437738 506128 437772
rect 506162 437738 506181 437772
rect 505711 437704 505730 437738
rect 505764 437722 506181 437738
rect 505764 437704 505877 437722
rect 505711 437688 505877 437704
rect 505911 437688 505978 437722
rect 506012 437688 506181 437722
rect 505711 437682 506181 437688
rect 505711 437648 506128 437682
rect 506162 437648 506181 437682
rect 505711 437614 505730 437648
rect 505764 437632 506181 437648
rect 505764 437614 505877 437632
rect 505711 437598 505877 437614
rect 505911 437598 505978 437632
rect 506012 437598 506181 437632
rect 505711 437592 506181 437598
rect 505711 437558 506128 437592
rect 506162 437558 506181 437592
rect 505711 437524 505730 437558
rect 505764 437542 506181 437558
rect 505764 437524 505877 437542
rect 505711 437508 505877 437524
rect 505911 437508 505978 437542
rect 506012 437508 506181 437542
rect 505711 437502 506181 437508
rect 504423 437434 504442 437468
rect 504476 437452 504893 437468
rect 504476 437434 504589 437452
rect 504423 437429 504589 437434
rect 503436 437418 504589 437429
rect 504623 437418 504690 437452
rect 504724 437429 504893 437452
rect 505711 437468 506128 437502
rect 506162 437468 506181 437502
rect 506243 438124 506937 438185
rect 506243 438090 506304 438124
rect 506338 438112 506394 438124
rect 506428 438112 506484 438124
rect 506518 438112 506574 438124
rect 506350 438090 506394 438112
rect 506450 438090 506484 438112
rect 506550 438090 506574 438112
rect 506608 438112 506664 438124
rect 506608 438090 506616 438112
rect 506243 438078 506316 438090
rect 506350 438078 506416 438090
rect 506450 438078 506516 438090
rect 506550 438078 506616 438090
rect 506650 438090 506664 438112
rect 506698 438112 506754 438124
rect 506698 438090 506716 438112
rect 506650 438078 506716 438090
rect 506750 438090 506754 438112
rect 506788 438112 506844 438124
rect 506788 438090 506816 438112
rect 506878 438090 506937 438124
rect 506750 438078 506816 438090
rect 506850 438078 506937 438090
rect 506243 438034 506937 438078
rect 506243 438000 506304 438034
rect 506338 438012 506394 438034
rect 506428 438012 506484 438034
rect 506518 438012 506574 438034
rect 506350 438000 506394 438012
rect 506450 438000 506484 438012
rect 506550 438000 506574 438012
rect 506608 438012 506664 438034
rect 506608 438000 506616 438012
rect 506243 437978 506316 438000
rect 506350 437978 506416 438000
rect 506450 437978 506516 438000
rect 506550 437978 506616 438000
rect 506650 438000 506664 438012
rect 506698 438012 506754 438034
rect 506698 438000 506716 438012
rect 506650 437978 506716 438000
rect 506750 438000 506754 438012
rect 506788 438012 506844 438034
rect 506788 438000 506816 438012
rect 506878 438000 506937 438034
rect 506750 437978 506816 438000
rect 506850 437978 506937 438000
rect 506243 437944 506937 437978
rect 506243 437910 506304 437944
rect 506338 437912 506394 437944
rect 506428 437912 506484 437944
rect 506518 437912 506574 437944
rect 506350 437910 506394 437912
rect 506450 437910 506484 437912
rect 506550 437910 506574 437912
rect 506608 437912 506664 437944
rect 506608 437910 506616 437912
rect 506243 437878 506316 437910
rect 506350 437878 506416 437910
rect 506450 437878 506516 437910
rect 506550 437878 506616 437910
rect 506650 437910 506664 437912
rect 506698 437912 506754 437944
rect 506698 437910 506716 437912
rect 506650 437878 506716 437910
rect 506750 437910 506754 437912
rect 506788 437912 506844 437944
rect 506788 437910 506816 437912
rect 506878 437910 506937 437944
rect 506750 437878 506816 437910
rect 506850 437878 506937 437910
rect 506243 437854 506937 437878
rect 506243 437820 506304 437854
rect 506338 437820 506394 437854
rect 506428 437820 506484 437854
rect 506518 437820 506574 437854
rect 506608 437820 506664 437854
rect 506698 437820 506754 437854
rect 506788 437820 506844 437854
rect 506878 437820 506937 437854
rect 506243 437812 506937 437820
rect 506243 437778 506316 437812
rect 506350 437778 506416 437812
rect 506450 437778 506516 437812
rect 506550 437778 506616 437812
rect 506650 437778 506716 437812
rect 506750 437778 506816 437812
rect 506850 437778 506937 437812
rect 506243 437764 506937 437778
rect 506243 437730 506304 437764
rect 506338 437730 506394 437764
rect 506428 437730 506484 437764
rect 506518 437730 506574 437764
rect 506608 437730 506664 437764
rect 506698 437730 506754 437764
rect 506788 437730 506844 437764
rect 506878 437730 506937 437764
rect 506243 437712 506937 437730
rect 506243 437678 506316 437712
rect 506350 437678 506416 437712
rect 506450 437678 506516 437712
rect 506550 437678 506616 437712
rect 506650 437678 506716 437712
rect 506750 437678 506816 437712
rect 506850 437678 506937 437712
rect 506243 437674 506937 437678
rect 506243 437640 506304 437674
rect 506338 437640 506394 437674
rect 506428 437640 506484 437674
rect 506518 437640 506574 437674
rect 506608 437640 506664 437674
rect 506698 437640 506754 437674
rect 506788 437640 506844 437674
rect 506878 437640 506937 437674
rect 506243 437612 506937 437640
rect 506243 437584 506316 437612
rect 506350 437584 506416 437612
rect 506450 437584 506516 437612
rect 506550 437584 506616 437612
rect 506243 437550 506304 437584
rect 506350 437578 506394 437584
rect 506450 437578 506484 437584
rect 506550 437578 506574 437584
rect 506338 437550 506394 437578
rect 506428 437550 506484 437578
rect 506518 437550 506574 437578
rect 506608 437578 506616 437584
rect 506650 437584 506716 437612
rect 506650 437578 506664 437584
rect 506608 437550 506664 437578
rect 506698 437578 506716 437584
rect 506750 437584 506816 437612
rect 506850 437584 506937 437612
rect 506750 437578 506754 437584
rect 506698 437550 506754 437578
rect 506788 437578 506816 437584
rect 506788 437550 506844 437578
rect 506878 437550 506937 437584
rect 506243 437491 506937 437550
rect 506999 438154 507018 438188
rect 507052 438172 507469 438188
rect 508287 438228 508453 438247
rect 508487 438228 508554 438262
rect 508588 438247 509741 438262
rect 508588 438228 508757 438247
rect 508287 438222 508757 438228
rect 508287 438188 508704 438222
rect 508738 438188 508757 438222
rect 507052 438154 507165 438172
rect 506999 438138 507165 438154
rect 507199 438138 507266 438172
rect 507300 438138 507469 438172
rect 506999 438132 507469 438138
rect 506999 438098 507416 438132
rect 507450 438098 507469 438132
rect 506999 438064 507018 438098
rect 507052 438082 507469 438098
rect 507052 438064 507165 438082
rect 506999 438048 507165 438064
rect 507199 438048 507266 438082
rect 507300 438048 507469 438082
rect 506999 438042 507469 438048
rect 506999 438008 507416 438042
rect 507450 438008 507469 438042
rect 506999 437974 507018 438008
rect 507052 437992 507469 438008
rect 507052 437974 507165 437992
rect 506999 437958 507165 437974
rect 507199 437958 507266 437992
rect 507300 437958 507469 437992
rect 506999 437952 507469 437958
rect 506999 437918 507416 437952
rect 507450 437918 507469 437952
rect 506999 437884 507018 437918
rect 507052 437902 507469 437918
rect 507052 437884 507165 437902
rect 506999 437868 507165 437884
rect 507199 437868 507266 437902
rect 507300 437868 507469 437902
rect 506999 437862 507469 437868
rect 506999 437828 507416 437862
rect 507450 437828 507469 437862
rect 506999 437794 507018 437828
rect 507052 437812 507469 437828
rect 507052 437794 507165 437812
rect 506999 437778 507165 437794
rect 507199 437778 507266 437812
rect 507300 437778 507469 437812
rect 506999 437772 507469 437778
rect 506999 437738 507416 437772
rect 507450 437738 507469 437772
rect 506999 437704 507018 437738
rect 507052 437722 507469 437738
rect 507052 437704 507165 437722
rect 506999 437688 507165 437704
rect 507199 437688 507266 437722
rect 507300 437688 507469 437722
rect 506999 437682 507469 437688
rect 506999 437648 507416 437682
rect 507450 437648 507469 437682
rect 506999 437614 507018 437648
rect 507052 437632 507469 437648
rect 507052 437614 507165 437632
rect 506999 437598 507165 437614
rect 507199 437598 507266 437632
rect 507300 437598 507469 437632
rect 506999 437592 507469 437598
rect 506999 437558 507416 437592
rect 507450 437558 507469 437592
rect 506999 437524 507018 437558
rect 507052 437542 507469 437558
rect 507052 437524 507165 437542
rect 506999 437508 507165 437524
rect 507199 437508 507266 437542
rect 507300 437508 507469 437542
rect 506999 437502 507469 437508
rect 505711 437434 505730 437468
rect 505764 437452 506181 437468
rect 505764 437434 505877 437452
rect 505711 437429 505877 437434
rect 504724 437418 505877 437429
rect 505911 437418 505978 437452
rect 506012 437429 506181 437452
rect 506999 437468 507416 437502
rect 507450 437468 507469 437502
rect 507531 438124 508225 438185
rect 507531 438090 507592 438124
rect 507626 438112 507682 438124
rect 507716 438112 507772 438124
rect 507806 438112 507862 438124
rect 507638 438090 507682 438112
rect 507738 438090 507772 438112
rect 507838 438090 507862 438112
rect 507896 438112 507952 438124
rect 507896 438090 507904 438112
rect 507531 438078 507604 438090
rect 507638 438078 507704 438090
rect 507738 438078 507804 438090
rect 507838 438078 507904 438090
rect 507938 438090 507952 438112
rect 507986 438112 508042 438124
rect 507986 438090 508004 438112
rect 507938 438078 508004 438090
rect 508038 438090 508042 438112
rect 508076 438112 508132 438124
rect 508076 438090 508104 438112
rect 508166 438090 508225 438124
rect 508038 438078 508104 438090
rect 508138 438078 508225 438090
rect 507531 438034 508225 438078
rect 507531 438000 507592 438034
rect 507626 438012 507682 438034
rect 507716 438012 507772 438034
rect 507806 438012 507862 438034
rect 507638 438000 507682 438012
rect 507738 438000 507772 438012
rect 507838 438000 507862 438012
rect 507896 438012 507952 438034
rect 507896 438000 507904 438012
rect 507531 437978 507604 438000
rect 507638 437978 507704 438000
rect 507738 437978 507804 438000
rect 507838 437978 507904 438000
rect 507938 438000 507952 438012
rect 507986 438012 508042 438034
rect 507986 438000 508004 438012
rect 507938 437978 508004 438000
rect 508038 438000 508042 438012
rect 508076 438012 508132 438034
rect 508076 438000 508104 438012
rect 508166 438000 508225 438034
rect 508038 437978 508104 438000
rect 508138 437978 508225 438000
rect 507531 437944 508225 437978
rect 507531 437910 507592 437944
rect 507626 437912 507682 437944
rect 507716 437912 507772 437944
rect 507806 437912 507862 437944
rect 507638 437910 507682 437912
rect 507738 437910 507772 437912
rect 507838 437910 507862 437912
rect 507896 437912 507952 437944
rect 507896 437910 507904 437912
rect 507531 437878 507604 437910
rect 507638 437878 507704 437910
rect 507738 437878 507804 437910
rect 507838 437878 507904 437910
rect 507938 437910 507952 437912
rect 507986 437912 508042 437944
rect 507986 437910 508004 437912
rect 507938 437878 508004 437910
rect 508038 437910 508042 437912
rect 508076 437912 508132 437944
rect 508076 437910 508104 437912
rect 508166 437910 508225 437944
rect 508038 437878 508104 437910
rect 508138 437878 508225 437910
rect 507531 437854 508225 437878
rect 507531 437820 507592 437854
rect 507626 437820 507682 437854
rect 507716 437820 507772 437854
rect 507806 437820 507862 437854
rect 507896 437820 507952 437854
rect 507986 437820 508042 437854
rect 508076 437820 508132 437854
rect 508166 437820 508225 437854
rect 507531 437812 508225 437820
rect 507531 437778 507604 437812
rect 507638 437778 507704 437812
rect 507738 437778 507804 437812
rect 507838 437778 507904 437812
rect 507938 437778 508004 437812
rect 508038 437778 508104 437812
rect 508138 437778 508225 437812
rect 507531 437764 508225 437778
rect 507531 437730 507592 437764
rect 507626 437730 507682 437764
rect 507716 437730 507772 437764
rect 507806 437730 507862 437764
rect 507896 437730 507952 437764
rect 507986 437730 508042 437764
rect 508076 437730 508132 437764
rect 508166 437730 508225 437764
rect 507531 437712 508225 437730
rect 507531 437678 507604 437712
rect 507638 437678 507704 437712
rect 507738 437678 507804 437712
rect 507838 437678 507904 437712
rect 507938 437678 508004 437712
rect 508038 437678 508104 437712
rect 508138 437678 508225 437712
rect 507531 437674 508225 437678
rect 507531 437640 507592 437674
rect 507626 437640 507682 437674
rect 507716 437640 507772 437674
rect 507806 437640 507862 437674
rect 507896 437640 507952 437674
rect 507986 437640 508042 437674
rect 508076 437640 508132 437674
rect 508166 437640 508225 437674
rect 507531 437612 508225 437640
rect 507531 437584 507604 437612
rect 507638 437584 507704 437612
rect 507738 437584 507804 437612
rect 507838 437584 507904 437612
rect 507531 437550 507592 437584
rect 507638 437578 507682 437584
rect 507738 437578 507772 437584
rect 507838 437578 507862 437584
rect 507626 437550 507682 437578
rect 507716 437550 507772 437578
rect 507806 437550 507862 437578
rect 507896 437578 507904 437584
rect 507938 437584 508004 437612
rect 507938 437578 507952 437584
rect 507896 437550 507952 437578
rect 507986 437578 508004 437584
rect 508038 437584 508104 437612
rect 508138 437584 508225 437612
rect 508038 437578 508042 437584
rect 507986 437550 508042 437578
rect 508076 437578 508104 437584
rect 508076 437550 508132 437578
rect 508166 437550 508225 437584
rect 507531 437491 508225 437550
rect 508287 438154 508306 438188
rect 508340 438172 508757 438188
rect 509575 438228 509741 438247
rect 509775 438228 509842 438262
rect 509876 438247 511029 438262
rect 509876 438228 510045 438247
rect 509575 438222 510045 438228
rect 509575 438188 509992 438222
rect 510026 438188 510045 438222
rect 508340 438154 508453 438172
rect 508287 438138 508453 438154
rect 508487 438138 508554 438172
rect 508588 438138 508757 438172
rect 508287 438132 508757 438138
rect 508287 438098 508704 438132
rect 508738 438098 508757 438132
rect 508287 438064 508306 438098
rect 508340 438082 508757 438098
rect 508340 438064 508453 438082
rect 508287 438048 508453 438064
rect 508487 438048 508554 438082
rect 508588 438048 508757 438082
rect 508287 438042 508757 438048
rect 508287 438008 508704 438042
rect 508738 438008 508757 438042
rect 508287 437974 508306 438008
rect 508340 437992 508757 438008
rect 508340 437974 508453 437992
rect 508287 437958 508453 437974
rect 508487 437958 508554 437992
rect 508588 437958 508757 437992
rect 508287 437952 508757 437958
rect 508287 437918 508704 437952
rect 508738 437918 508757 437952
rect 508287 437884 508306 437918
rect 508340 437902 508757 437918
rect 508340 437884 508453 437902
rect 508287 437868 508453 437884
rect 508487 437868 508554 437902
rect 508588 437868 508757 437902
rect 508287 437862 508757 437868
rect 508287 437828 508704 437862
rect 508738 437828 508757 437862
rect 508287 437794 508306 437828
rect 508340 437812 508757 437828
rect 508340 437794 508453 437812
rect 508287 437778 508453 437794
rect 508487 437778 508554 437812
rect 508588 437778 508757 437812
rect 508287 437772 508757 437778
rect 508287 437738 508704 437772
rect 508738 437738 508757 437772
rect 508287 437704 508306 437738
rect 508340 437722 508757 437738
rect 508340 437704 508453 437722
rect 508287 437688 508453 437704
rect 508487 437688 508554 437722
rect 508588 437688 508757 437722
rect 508287 437682 508757 437688
rect 508287 437648 508704 437682
rect 508738 437648 508757 437682
rect 508287 437614 508306 437648
rect 508340 437632 508757 437648
rect 508340 437614 508453 437632
rect 508287 437598 508453 437614
rect 508487 437598 508554 437632
rect 508588 437598 508757 437632
rect 508287 437592 508757 437598
rect 508287 437558 508704 437592
rect 508738 437558 508757 437592
rect 508287 437524 508306 437558
rect 508340 437542 508757 437558
rect 508340 437524 508453 437542
rect 508287 437508 508453 437524
rect 508487 437508 508554 437542
rect 508588 437508 508757 437542
rect 508287 437502 508757 437508
rect 506999 437434 507018 437468
rect 507052 437452 507469 437468
rect 507052 437434 507165 437452
rect 506999 437429 507165 437434
rect 506012 437418 507165 437429
rect 507199 437418 507266 437452
rect 507300 437429 507469 437452
rect 508287 437468 508704 437502
rect 508738 437468 508757 437502
rect 508819 438124 509513 438185
rect 508819 438090 508880 438124
rect 508914 438112 508970 438124
rect 509004 438112 509060 438124
rect 509094 438112 509150 438124
rect 508926 438090 508970 438112
rect 509026 438090 509060 438112
rect 509126 438090 509150 438112
rect 509184 438112 509240 438124
rect 509184 438090 509192 438112
rect 508819 438078 508892 438090
rect 508926 438078 508992 438090
rect 509026 438078 509092 438090
rect 509126 438078 509192 438090
rect 509226 438090 509240 438112
rect 509274 438112 509330 438124
rect 509274 438090 509292 438112
rect 509226 438078 509292 438090
rect 509326 438090 509330 438112
rect 509364 438112 509420 438124
rect 509364 438090 509392 438112
rect 509454 438090 509513 438124
rect 509326 438078 509392 438090
rect 509426 438078 509513 438090
rect 508819 438034 509513 438078
rect 508819 438000 508880 438034
rect 508914 438012 508970 438034
rect 509004 438012 509060 438034
rect 509094 438012 509150 438034
rect 508926 438000 508970 438012
rect 509026 438000 509060 438012
rect 509126 438000 509150 438012
rect 509184 438012 509240 438034
rect 509184 438000 509192 438012
rect 508819 437978 508892 438000
rect 508926 437978 508992 438000
rect 509026 437978 509092 438000
rect 509126 437978 509192 438000
rect 509226 438000 509240 438012
rect 509274 438012 509330 438034
rect 509274 438000 509292 438012
rect 509226 437978 509292 438000
rect 509326 438000 509330 438012
rect 509364 438012 509420 438034
rect 509364 438000 509392 438012
rect 509454 438000 509513 438034
rect 509326 437978 509392 438000
rect 509426 437978 509513 438000
rect 508819 437944 509513 437978
rect 508819 437910 508880 437944
rect 508914 437912 508970 437944
rect 509004 437912 509060 437944
rect 509094 437912 509150 437944
rect 508926 437910 508970 437912
rect 509026 437910 509060 437912
rect 509126 437910 509150 437912
rect 509184 437912 509240 437944
rect 509184 437910 509192 437912
rect 508819 437878 508892 437910
rect 508926 437878 508992 437910
rect 509026 437878 509092 437910
rect 509126 437878 509192 437910
rect 509226 437910 509240 437912
rect 509274 437912 509330 437944
rect 509274 437910 509292 437912
rect 509226 437878 509292 437910
rect 509326 437910 509330 437912
rect 509364 437912 509420 437944
rect 509364 437910 509392 437912
rect 509454 437910 509513 437944
rect 509326 437878 509392 437910
rect 509426 437878 509513 437910
rect 508819 437854 509513 437878
rect 508819 437820 508880 437854
rect 508914 437820 508970 437854
rect 509004 437820 509060 437854
rect 509094 437820 509150 437854
rect 509184 437820 509240 437854
rect 509274 437820 509330 437854
rect 509364 437820 509420 437854
rect 509454 437820 509513 437854
rect 508819 437812 509513 437820
rect 508819 437778 508892 437812
rect 508926 437778 508992 437812
rect 509026 437778 509092 437812
rect 509126 437778 509192 437812
rect 509226 437778 509292 437812
rect 509326 437778 509392 437812
rect 509426 437778 509513 437812
rect 508819 437764 509513 437778
rect 508819 437730 508880 437764
rect 508914 437730 508970 437764
rect 509004 437730 509060 437764
rect 509094 437730 509150 437764
rect 509184 437730 509240 437764
rect 509274 437730 509330 437764
rect 509364 437730 509420 437764
rect 509454 437730 509513 437764
rect 508819 437712 509513 437730
rect 508819 437678 508892 437712
rect 508926 437678 508992 437712
rect 509026 437678 509092 437712
rect 509126 437678 509192 437712
rect 509226 437678 509292 437712
rect 509326 437678 509392 437712
rect 509426 437678 509513 437712
rect 508819 437674 509513 437678
rect 508819 437640 508880 437674
rect 508914 437640 508970 437674
rect 509004 437640 509060 437674
rect 509094 437640 509150 437674
rect 509184 437640 509240 437674
rect 509274 437640 509330 437674
rect 509364 437640 509420 437674
rect 509454 437640 509513 437674
rect 508819 437612 509513 437640
rect 508819 437584 508892 437612
rect 508926 437584 508992 437612
rect 509026 437584 509092 437612
rect 509126 437584 509192 437612
rect 508819 437550 508880 437584
rect 508926 437578 508970 437584
rect 509026 437578 509060 437584
rect 509126 437578 509150 437584
rect 508914 437550 508970 437578
rect 509004 437550 509060 437578
rect 509094 437550 509150 437578
rect 509184 437578 509192 437584
rect 509226 437584 509292 437612
rect 509226 437578 509240 437584
rect 509184 437550 509240 437578
rect 509274 437578 509292 437584
rect 509326 437584 509392 437612
rect 509426 437584 509513 437612
rect 509326 437578 509330 437584
rect 509274 437550 509330 437578
rect 509364 437578 509392 437584
rect 509364 437550 509420 437578
rect 509454 437550 509513 437584
rect 508819 437491 509513 437550
rect 509575 438154 509594 438188
rect 509628 438172 510045 438188
rect 510863 438228 511029 438247
rect 511063 438228 511130 438262
rect 511164 438247 512317 438262
rect 511164 438228 511333 438247
rect 510863 438222 511333 438228
rect 510863 438188 511280 438222
rect 511314 438188 511333 438222
rect 509628 438154 509741 438172
rect 509575 438138 509741 438154
rect 509775 438138 509842 438172
rect 509876 438138 510045 438172
rect 509575 438132 510045 438138
rect 509575 438098 509992 438132
rect 510026 438098 510045 438132
rect 509575 438064 509594 438098
rect 509628 438082 510045 438098
rect 509628 438064 509741 438082
rect 509575 438048 509741 438064
rect 509775 438048 509842 438082
rect 509876 438048 510045 438082
rect 509575 438042 510045 438048
rect 509575 438008 509992 438042
rect 510026 438008 510045 438042
rect 509575 437974 509594 438008
rect 509628 437992 510045 438008
rect 509628 437974 509741 437992
rect 509575 437958 509741 437974
rect 509775 437958 509842 437992
rect 509876 437958 510045 437992
rect 509575 437952 510045 437958
rect 509575 437918 509992 437952
rect 510026 437918 510045 437952
rect 509575 437884 509594 437918
rect 509628 437902 510045 437918
rect 509628 437884 509741 437902
rect 509575 437868 509741 437884
rect 509775 437868 509842 437902
rect 509876 437868 510045 437902
rect 509575 437862 510045 437868
rect 509575 437828 509992 437862
rect 510026 437828 510045 437862
rect 509575 437794 509594 437828
rect 509628 437812 510045 437828
rect 509628 437794 509741 437812
rect 509575 437778 509741 437794
rect 509775 437778 509842 437812
rect 509876 437778 510045 437812
rect 509575 437772 510045 437778
rect 509575 437738 509992 437772
rect 510026 437738 510045 437772
rect 509575 437704 509594 437738
rect 509628 437722 510045 437738
rect 509628 437704 509741 437722
rect 509575 437688 509741 437704
rect 509775 437688 509842 437722
rect 509876 437688 510045 437722
rect 509575 437682 510045 437688
rect 509575 437648 509992 437682
rect 510026 437648 510045 437682
rect 509575 437614 509594 437648
rect 509628 437632 510045 437648
rect 509628 437614 509741 437632
rect 509575 437598 509741 437614
rect 509775 437598 509842 437632
rect 509876 437598 510045 437632
rect 509575 437592 510045 437598
rect 509575 437558 509992 437592
rect 510026 437558 510045 437592
rect 509575 437524 509594 437558
rect 509628 437542 510045 437558
rect 509628 437524 509741 437542
rect 509575 437508 509741 437524
rect 509775 437508 509842 437542
rect 509876 437508 510045 437542
rect 509575 437502 510045 437508
rect 508287 437434 508306 437468
rect 508340 437452 508757 437468
rect 508340 437434 508453 437452
rect 508287 437429 508453 437434
rect 507300 437418 508453 437429
rect 508487 437418 508554 437452
rect 508588 437429 508757 437452
rect 509575 437468 509992 437502
rect 510026 437468 510045 437502
rect 510107 438124 510801 438185
rect 510107 438090 510168 438124
rect 510202 438112 510258 438124
rect 510292 438112 510348 438124
rect 510382 438112 510438 438124
rect 510214 438090 510258 438112
rect 510314 438090 510348 438112
rect 510414 438090 510438 438112
rect 510472 438112 510528 438124
rect 510472 438090 510480 438112
rect 510107 438078 510180 438090
rect 510214 438078 510280 438090
rect 510314 438078 510380 438090
rect 510414 438078 510480 438090
rect 510514 438090 510528 438112
rect 510562 438112 510618 438124
rect 510562 438090 510580 438112
rect 510514 438078 510580 438090
rect 510614 438090 510618 438112
rect 510652 438112 510708 438124
rect 510652 438090 510680 438112
rect 510742 438090 510801 438124
rect 510614 438078 510680 438090
rect 510714 438078 510801 438090
rect 510107 438034 510801 438078
rect 510107 438000 510168 438034
rect 510202 438012 510258 438034
rect 510292 438012 510348 438034
rect 510382 438012 510438 438034
rect 510214 438000 510258 438012
rect 510314 438000 510348 438012
rect 510414 438000 510438 438012
rect 510472 438012 510528 438034
rect 510472 438000 510480 438012
rect 510107 437978 510180 438000
rect 510214 437978 510280 438000
rect 510314 437978 510380 438000
rect 510414 437978 510480 438000
rect 510514 438000 510528 438012
rect 510562 438012 510618 438034
rect 510562 438000 510580 438012
rect 510514 437978 510580 438000
rect 510614 438000 510618 438012
rect 510652 438012 510708 438034
rect 510652 438000 510680 438012
rect 510742 438000 510801 438034
rect 510614 437978 510680 438000
rect 510714 437978 510801 438000
rect 510107 437944 510801 437978
rect 510107 437910 510168 437944
rect 510202 437912 510258 437944
rect 510292 437912 510348 437944
rect 510382 437912 510438 437944
rect 510214 437910 510258 437912
rect 510314 437910 510348 437912
rect 510414 437910 510438 437912
rect 510472 437912 510528 437944
rect 510472 437910 510480 437912
rect 510107 437878 510180 437910
rect 510214 437878 510280 437910
rect 510314 437878 510380 437910
rect 510414 437878 510480 437910
rect 510514 437910 510528 437912
rect 510562 437912 510618 437944
rect 510562 437910 510580 437912
rect 510514 437878 510580 437910
rect 510614 437910 510618 437912
rect 510652 437912 510708 437944
rect 510652 437910 510680 437912
rect 510742 437910 510801 437944
rect 510614 437878 510680 437910
rect 510714 437878 510801 437910
rect 510107 437854 510801 437878
rect 510107 437820 510168 437854
rect 510202 437820 510258 437854
rect 510292 437820 510348 437854
rect 510382 437820 510438 437854
rect 510472 437820 510528 437854
rect 510562 437820 510618 437854
rect 510652 437820 510708 437854
rect 510742 437820 510801 437854
rect 510107 437812 510801 437820
rect 510107 437778 510180 437812
rect 510214 437778 510280 437812
rect 510314 437778 510380 437812
rect 510414 437778 510480 437812
rect 510514 437778 510580 437812
rect 510614 437778 510680 437812
rect 510714 437778 510801 437812
rect 510107 437764 510801 437778
rect 510107 437730 510168 437764
rect 510202 437730 510258 437764
rect 510292 437730 510348 437764
rect 510382 437730 510438 437764
rect 510472 437730 510528 437764
rect 510562 437730 510618 437764
rect 510652 437730 510708 437764
rect 510742 437730 510801 437764
rect 510107 437712 510801 437730
rect 510107 437678 510180 437712
rect 510214 437678 510280 437712
rect 510314 437678 510380 437712
rect 510414 437678 510480 437712
rect 510514 437678 510580 437712
rect 510614 437678 510680 437712
rect 510714 437678 510801 437712
rect 510107 437674 510801 437678
rect 510107 437640 510168 437674
rect 510202 437640 510258 437674
rect 510292 437640 510348 437674
rect 510382 437640 510438 437674
rect 510472 437640 510528 437674
rect 510562 437640 510618 437674
rect 510652 437640 510708 437674
rect 510742 437640 510801 437674
rect 510107 437612 510801 437640
rect 510107 437584 510180 437612
rect 510214 437584 510280 437612
rect 510314 437584 510380 437612
rect 510414 437584 510480 437612
rect 510107 437550 510168 437584
rect 510214 437578 510258 437584
rect 510314 437578 510348 437584
rect 510414 437578 510438 437584
rect 510202 437550 510258 437578
rect 510292 437550 510348 437578
rect 510382 437550 510438 437578
rect 510472 437578 510480 437584
rect 510514 437584 510580 437612
rect 510514 437578 510528 437584
rect 510472 437550 510528 437578
rect 510562 437578 510580 437584
rect 510614 437584 510680 437612
rect 510714 437584 510801 437612
rect 510614 437578 510618 437584
rect 510562 437550 510618 437578
rect 510652 437578 510680 437584
rect 510652 437550 510708 437578
rect 510742 437550 510801 437584
rect 510107 437491 510801 437550
rect 510863 438154 510882 438188
rect 510916 438172 511333 438188
rect 512151 438228 512317 438247
rect 512351 438228 512418 438262
rect 512452 438247 513605 438262
rect 512452 438228 512621 438247
rect 512151 438222 512621 438228
rect 512151 438188 512568 438222
rect 512602 438188 512621 438222
rect 510916 438154 511029 438172
rect 510863 438138 511029 438154
rect 511063 438138 511130 438172
rect 511164 438138 511333 438172
rect 510863 438132 511333 438138
rect 510863 438098 511280 438132
rect 511314 438098 511333 438132
rect 510863 438064 510882 438098
rect 510916 438082 511333 438098
rect 510916 438064 511029 438082
rect 510863 438048 511029 438064
rect 511063 438048 511130 438082
rect 511164 438048 511333 438082
rect 510863 438042 511333 438048
rect 510863 438008 511280 438042
rect 511314 438008 511333 438042
rect 510863 437974 510882 438008
rect 510916 437992 511333 438008
rect 510916 437974 511029 437992
rect 510863 437958 511029 437974
rect 511063 437958 511130 437992
rect 511164 437958 511333 437992
rect 510863 437952 511333 437958
rect 510863 437918 511280 437952
rect 511314 437918 511333 437952
rect 510863 437884 510882 437918
rect 510916 437902 511333 437918
rect 510916 437884 511029 437902
rect 510863 437868 511029 437884
rect 511063 437868 511130 437902
rect 511164 437868 511333 437902
rect 510863 437862 511333 437868
rect 510863 437828 511280 437862
rect 511314 437828 511333 437862
rect 510863 437794 510882 437828
rect 510916 437812 511333 437828
rect 510916 437794 511029 437812
rect 510863 437778 511029 437794
rect 511063 437778 511130 437812
rect 511164 437778 511333 437812
rect 510863 437772 511333 437778
rect 510863 437738 511280 437772
rect 511314 437738 511333 437772
rect 510863 437704 510882 437738
rect 510916 437722 511333 437738
rect 510916 437704 511029 437722
rect 510863 437688 511029 437704
rect 511063 437688 511130 437722
rect 511164 437688 511333 437722
rect 510863 437682 511333 437688
rect 510863 437648 511280 437682
rect 511314 437648 511333 437682
rect 510863 437614 510882 437648
rect 510916 437632 511333 437648
rect 510916 437614 511029 437632
rect 510863 437598 511029 437614
rect 511063 437598 511130 437632
rect 511164 437598 511333 437632
rect 510863 437592 511333 437598
rect 510863 437558 511280 437592
rect 511314 437558 511333 437592
rect 510863 437524 510882 437558
rect 510916 437542 511333 437558
rect 510916 437524 511029 437542
rect 510863 437508 511029 437524
rect 511063 437508 511130 437542
rect 511164 437508 511333 437542
rect 510863 437502 511333 437508
rect 509575 437434 509594 437468
rect 509628 437452 510045 437468
rect 509628 437434 509741 437452
rect 509575 437429 509741 437434
rect 508588 437418 509741 437429
rect 509775 437418 509842 437452
rect 509876 437429 510045 437452
rect 510863 437468 511280 437502
rect 511314 437468 511333 437502
rect 511395 438124 512089 438185
rect 511395 438090 511456 438124
rect 511490 438112 511546 438124
rect 511580 438112 511636 438124
rect 511670 438112 511726 438124
rect 511502 438090 511546 438112
rect 511602 438090 511636 438112
rect 511702 438090 511726 438112
rect 511760 438112 511816 438124
rect 511760 438090 511768 438112
rect 511395 438078 511468 438090
rect 511502 438078 511568 438090
rect 511602 438078 511668 438090
rect 511702 438078 511768 438090
rect 511802 438090 511816 438112
rect 511850 438112 511906 438124
rect 511850 438090 511868 438112
rect 511802 438078 511868 438090
rect 511902 438090 511906 438112
rect 511940 438112 511996 438124
rect 511940 438090 511968 438112
rect 512030 438090 512089 438124
rect 511902 438078 511968 438090
rect 512002 438078 512089 438090
rect 511395 438034 512089 438078
rect 511395 438000 511456 438034
rect 511490 438012 511546 438034
rect 511580 438012 511636 438034
rect 511670 438012 511726 438034
rect 511502 438000 511546 438012
rect 511602 438000 511636 438012
rect 511702 438000 511726 438012
rect 511760 438012 511816 438034
rect 511760 438000 511768 438012
rect 511395 437978 511468 438000
rect 511502 437978 511568 438000
rect 511602 437978 511668 438000
rect 511702 437978 511768 438000
rect 511802 438000 511816 438012
rect 511850 438012 511906 438034
rect 511850 438000 511868 438012
rect 511802 437978 511868 438000
rect 511902 438000 511906 438012
rect 511940 438012 511996 438034
rect 511940 438000 511968 438012
rect 512030 438000 512089 438034
rect 511902 437978 511968 438000
rect 512002 437978 512089 438000
rect 511395 437944 512089 437978
rect 511395 437910 511456 437944
rect 511490 437912 511546 437944
rect 511580 437912 511636 437944
rect 511670 437912 511726 437944
rect 511502 437910 511546 437912
rect 511602 437910 511636 437912
rect 511702 437910 511726 437912
rect 511760 437912 511816 437944
rect 511760 437910 511768 437912
rect 511395 437878 511468 437910
rect 511502 437878 511568 437910
rect 511602 437878 511668 437910
rect 511702 437878 511768 437910
rect 511802 437910 511816 437912
rect 511850 437912 511906 437944
rect 511850 437910 511868 437912
rect 511802 437878 511868 437910
rect 511902 437910 511906 437912
rect 511940 437912 511996 437944
rect 511940 437910 511968 437912
rect 512030 437910 512089 437944
rect 511902 437878 511968 437910
rect 512002 437878 512089 437910
rect 511395 437854 512089 437878
rect 511395 437820 511456 437854
rect 511490 437820 511546 437854
rect 511580 437820 511636 437854
rect 511670 437820 511726 437854
rect 511760 437820 511816 437854
rect 511850 437820 511906 437854
rect 511940 437820 511996 437854
rect 512030 437820 512089 437854
rect 511395 437812 512089 437820
rect 511395 437778 511468 437812
rect 511502 437778 511568 437812
rect 511602 437778 511668 437812
rect 511702 437778 511768 437812
rect 511802 437778 511868 437812
rect 511902 437778 511968 437812
rect 512002 437778 512089 437812
rect 511395 437764 512089 437778
rect 511395 437730 511456 437764
rect 511490 437730 511546 437764
rect 511580 437730 511636 437764
rect 511670 437730 511726 437764
rect 511760 437730 511816 437764
rect 511850 437730 511906 437764
rect 511940 437730 511996 437764
rect 512030 437730 512089 437764
rect 511395 437712 512089 437730
rect 511395 437678 511468 437712
rect 511502 437678 511568 437712
rect 511602 437678 511668 437712
rect 511702 437678 511768 437712
rect 511802 437678 511868 437712
rect 511902 437678 511968 437712
rect 512002 437678 512089 437712
rect 511395 437674 512089 437678
rect 511395 437640 511456 437674
rect 511490 437640 511546 437674
rect 511580 437640 511636 437674
rect 511670 437640 511726 437674
rect 511760 437640 511816 437674
rect 511850 437640 511906 437674
rect 511940 437640 511996 437674
rect 512030 437640 512089 437674
rect 511395 437612 512089 437640
rect 511395 437584 511468 437612
rect 511502 437584 511568 437612
rect 511602 437584 511668 437612
rect 511702 437584 511768 437612
rect 511395 437550 511456 437584
rect 511502 437578 511546 437584
rect 511602 437578 511636 437584
rect 511702 437578 511726 437584
rect 511490 437550 511546 437578
rect 511580 437550 511636 437578
rect 511670 437550 511726 437578
rect 511760 437578 511768 437584
rect 511802 437584 511868 437612
rect 511802 437578 511816 437584
rect 511760 437550 511816 437578
rect 511850 437578 511868 437584
rect 511902 437584 511968 437612
rect 512002 437584 512089 437612
rect 511902 437578 511906 437584
rect 511850 437550 511906 437578
rect 511940 437578 511968 437584
rect 511940 437550 511996 437578
rect 512030 437550 512089 437584
rect 511395 437491 512089 437550
rect 512151 438154 512170 438188
rect 512204 438172 512621 438188
rect 513439 438228 513605 438247
rect 513639 438228 513674 438262
rect 513439 438188 513674 438228
rect 512204 438154 512317 438172
rect 512151 438138 512317 438154
rect 512351 438138 512418 438172
rect 512452 438138 512621 438172
rect 512151 438132 512621 438138
rect 512151 438098 512568 438132
rect 512602 438098 512621 438132
rect 512151 438064 512170 438098
rect 512204 438082 512621 438098
rect 512204 438064 512317 438082
rect 512151 438048 512317 438064
rect 512351 438048 512418 438082
rect 512452 438048 512621 438082
rect 512151 438042 512621 438048
rect 512151 438008 512568 438042
rect 512602 438008 512621 438042
rect 512151 437974 512170 438008
rect 512204 437992 512621 438008
rect 512204 437974 512317 437992
rect 512151 437958 512317 437974
rect 512351 437958 512418 437992
rect 512452 437958 512621 437992
rect 512151 437952 512621 437958
rect 512151 437918 512568 437952
rect 512602 437918 512621 437952
rect 512151 437884 512170 437918
rect 512204 437902 512621 437918
rect 512204 437884 512317 437902
rect 512151 437868 512317 437884
rect 512351 437868 512418 437902
rect 512452 437868 512621 437902
rect 512151 437862 512621 437868
rect 512151 437828 512568 437862
rect 512602 437828 512621 437862
rect 512151 437794 512170 437828
rect 512204 437812 512621 437828
rect 512204 437794 512317 437812
rect 512151 437778 512317 437794
rect 512351 437778 512418 437812
rect 512452 437778 512621 437812
rect 512151 437772 512621 437778
rect 512151 437738 512568 437772
rect 512602 437738 512621 437772
rect 512151 437704 512170 437738
rect 512204 437722 512621 437738
rect 512204 437704 512317 437722
rect 512151 437688 512317 437704
rect 512351 437688 512418 437722
rect 512452 437688 512621 437722
rect 512151 437682 512621 437688
rect 512151 437648 512568 437682
rect 512602 437648 512621 437682
rect 512151 437614 512170 437648
rect 512204 437632 512621 437648
rect 512204 437614 512317 437632
rect 512151 437598 512317 437614
rect 512351 437598 512418 437632
rect 512452 437598 512621 437632
rect 512151 437592 512621 437598
rect 512151 437558 512568 437592
rect 512602 437558 512621 437592
rect 512151 437524 512170 437558
rect 512204 437542 512621 437558
rect 512204 437524 512317 437542
rect 512151 437508 512317 437524
rect 512351 437508 512418 437542
rect 512452 437508 512621 437542
rect 512151 437502 512621 437508
rect 510863 437434 510882 437468
rect 510916 437452 511333 437468
rect 510916 437434 511029 437452
rect 510863 437429 511029 437434
rect 509876 437418 511029 437429
rect 511063 437418 511130 437452
rect 511164 437429 511333 437452
rect 512151 437468 512568 437502
rect 512602 437468 512621 437502
rect 512683 438124 513377 438185
rect 512683 438090 512744 438124
rect 512778 438112 512834 438124
rect 512868 438112 512924 438124
rect 512958 438112 513014 438124
rect 512790 438090 512834 438112
rect 512890 438090 512924 438112
rect 512990 438090 513014 438112
rect 513048 438112 513104 438124
rect 513048 438090 513056 438112
rect 512683 438078 512756 438090
rect 512790 438078 512856 438090
rect 512890 438078 512956 438090
rect 512990 438078 513056 438090
rect 513090 438090 513104 438112
rect 513138 438112 513194 438124
rect 513138 438090 513156 438112
rect 513090 438078 513156 438090
rect 513190 438090 513194 438112
rect 513228 438112 513284 438124
rect 513228 438090 513256 438112
rect 513318 438090 513377 438124
rect 513190 438078 513256 438090
rect 513290 438078 513377 438090
rect 512683 438034 513377 438078
rect 512683 438000 512744 438034
rect 512778 438012 512834 438034
rect 512868 438012 512924 438034
rect 512958 438012 513014 438034
rect 512790 438000 512834 438012
rect 512890 438000 512924 438012
rect 512990 438000 513014 438012
rect 513048 438012 513104 438034
rect 513048 438000 513056 438012
rect 512683 437978 512756 438000
rect 512790 437978 512856 438000
rect 512890 437978 512956 438000
rect 512990 437978 513056 438000
rect 513090 438000 513104 438012
rect 513138 438012 513194 438034
rect 513138 438000 513156 438012
rect 513090 437978 513156 438000
rect 513190 438000 513194 438012
rect 513228 438012 513284 438034
rect 513228 438000 513256 438012
rect 513318 438000 513377 438034
rect 513190 437978 513256 438000
rect 513290 437978 513377 438000
rect 512683 437944 513377 437978
rect 512683 437910 512744 437944
rect 512778 437912 512834 437944
rect 512868 437912 512924 437944
rect 512958 437912 513014 437944
rect 512790 437910 512834 437912
rect 512890 437910 512924 437912
rect 512990 437910 513014 437912
rect 513048 437912 513104 437944
rect 513048 437910 513056 437912
rect 512683 437878 512756 437910
rect 512790 437878 512856 437910
rect 512890 437878 512956 437910
rect 512990 437878 513056 437910
rect 513090 437910 513104 437912
rect 513138 437912 513194 437944
rect 513138 437910 513156 437912
rect 513090 437878 513156 437910
rect 513190 437910 513194 437912
rect 513228 437912 513284 437944
rect 513228 437910 513256 437912
rect 513318 437910 513377 437944
rect 513190 437878 513256 437910
rect 513290 437878 513377 437910
rect 512683 437854 513377 437878
rect 512683 437820 512744 437854
rect 512778 437820 512834 437854
rect 512868 437820 512924 437854
rect 512958 437820 513014 437854
rect 513048 437820 513104 437854
rect 513138 437820 513194 437854
rect 513228 437820 513284 437854
rect 513318 437820 513377 437854
rect 512683 437812 513377 437820
rect 512683 437778 512756 437812
rect 512790 437778 512856 437812
rect 512890 437778 512956 437812
rect 512990 437778 513056 437812
rect 513090 437778 513156 437812
rect 513190 437778 513256 437812
rect 513290 437778 513377 437812
rect 512683 437764 513377 437778
rect 512683 437730 512744 437764
rect 512778 437730 512834 437764
rect 512868 437730 512924 437764
rect 512958 437730 513014 437764
rect 513048 437730 513104 437764
rect 513138 437730 513194 437764
rect 513228 437730 513284 437764
rect 513318 437730 513377 437764
rect 512683 437712 513377 437730
rect 512683 437678 512756 437712
rect 512790 437678 512856 437712
rect 512890 437678 512956 437712
rect 512990 437678 513056 437712
rect 513090 437678 513156 437712
rect 513190 437678 513256 437712
rect 513290 437678 513377 437712
rect 512683 437674 513377 437678
rect 512683 437640 512744 437674
rect 512778 437640 512834 437674
rect 512868 437640 512924 437674
rect 512958 437640 513014 437674
rect 513048 437640 513104 437674
rect 513138 437640 513194 437674
rect 513228 437640 513284 437674
rect 513318 437640 513377 437674
rect 512683 437612 513377 437640
rect 512683 437584 512756 437612
rect 512790 437584 512856 437612
rect 512890 437584 512956 437612
rect 512990 437584 513056 437612
rect 512683 437550 512744 437584
rect 512790 437578 512834 437584
rect 512890 437578 512924 437584
rect 512990 437578 513014 437584
rect 512778 437550 512834 437578
rect 512868 437550 512924 437578
rect 512958 437550 513014 437578
rect 513048 437578 513056 437584
rect 513090 437584 513156 437612
rect 513090 437578 513104 437584
rect 513048 437550 513104 437578
rect 513138 437578 513156 437584
rect 513190 437584 513256 437612
rect 513290 437584 513377 437612
rect 513190 437578 513194 437584
rect 513138 437550 513194 437578
rect 513228 437578 513256 437584
rect 513228 437550 513284 437578
rect 513318 437550 513377 437584
rect 512683 437491 513377 437550
rect 513439 438154 513458 438188
rect 513492 438172 513674 438188
rect 513492 438154 513605 438172
rect 513439 438138 513605 438154
rect 513639 438138 513674 438172
rect 513439 438098 513674 438138
rect 513439 438064 513458 438098
rect 513492 438082 513674 438098
rect 513492 438064 513605 438082
rect 513439 438048 513605 438064
rect 513639 438048 513674 438082
rect 513439 438008 513674 438048
rect 513439 437974 513458 438008
rect 513492 437992 513674 438008
rect 513492 437974 513605 437992
rect 513439 437958 513605 437974
rect 513639 437958 513674 437992
rect 513439 437918 513674 437958
rect 513439 437884 513458 437918
rect 513492 437902 513674 437918
rect 513492 437884 513605 437902
rect 513439 437868 513605 437884
rect 513639 437868 513674 437902
rect 513439 437828 513674 437868
rect 513439 437794 513458 437828
rect 513492 437812 513674 437828
rect 513492 437794 513605 437812
rect 513439 437778 513605 437794
rect 513639 437778 513674 437812
rect 513439 437738 513674 437778
rect 513439 437704 513458 437738
rect 513492 437722 513674 437738
rect 513492 437704 513605 437722
rect 513439 437688 513605 437704
rect 513639 437688 513674 437722
rect 513439 437648 513674 437688
rect 513439 437614 513458 437648
rect 513492 437632 513674 437648
rect 513492 437614 513605 437632
rect 513439 437598 513605 437614
rect 513639 437598 513674 437632
rect 513439 437558 513674 437598
rect 513439 437524 513458 437558
rect 513492 437542 513674 437558
rect 513492 437524 513605 437542
rect 513439 437508 513605 437524
rect 513639 437508 513674 437542
rect 512151 437434 512170 437468
rect 512204 437452 512621 437468
rect 512204 437434 512317 437452
rect 512151 437429 512317 437434
rect 511164 437418 512317 437429
rect 512351 437418 512418 437452
rect 512452 437429 512621 437452
rect 513439 437468 513674 437508
rect 513439 437434 513458 437468
rect 513492 437452 513674 437468
rect 513492 437434 513605 437452
rect 513439 437429 513605 437434
rect 512452 437418 513605 437429
rect 513639 437418 513674 437452
rect 503370 437410 513674 437418
rect 503370 437376 503646 437410
rect 503680 437376 503736 437410
rect 503770 437376 503826 437410
rect 503860 437376 503916 437410
rect 503950 437376 504006 437410
rect 504040 437376 504096 437410
rect 504130 437376 504186 437410
rect 504220 437376 504276 437410
rect 504310 437376 504366 437410
rect 504400 437376 504934 437410
rect 504968 437376 505024 437410
rect 505058 437376 505114 437410
rect 505148 437376 505204 437410
rect 505238 437376 505294 437410
rect 505328 437376 505384 437410
rect 505418 437376 505474 437410
rect 505508 437376 505564 437410
rect 505598 437376 505654 437410
rect 505688 437376 506222 437410
rect 506256 437376 506312 437410
rect 506346 437376 506402 437410
rect 506436 437376 506492 437410
rect 506526 437376 506582 437410
rect 506616 437376 506672 437410
rect 506706 437376 506762 437410
rect 506796 437376 506852 437410
rect 506886 437376 506942 437410
rect 506976 437376 507510 437410
rect 507544 437376 507600 437410
rect 507634 437376 507690 437410
rect 507724 437376 507780 437410
rect 507814 437376 507870 437410
rect 507904 437376 507960 437410
rect 507994 437376 508050 437410
rect 508084 437376 508140 437410
rect 508174 437376 508230 437410
rect 508264 437376 508798 437410
rect 508832 437376 508888 437410
rect 508922 437376 508978 437410
rect 509012 437376 509068 437410
rect 509102 437376 509158 437410
rect 509192 437376 509248 437410
rect 509282 437376 509338 437410
rect 509372 437376 509428 437410
rect 509462 437376 509518 437410
rect 509552 437376 510086 437410
rect 510120 437376 510176 437410
rect 510210 437376 510266 437410
rect 510300 437376 510356 437410
rect 510390 437376 510446 437410
rect 510480 437376 510536 437410
rect 510570 437376 510626 437410
rect 510660 437376 510716 437410
rect 510750 437376 510806 437410
rect 510840 437376 511374 437410
rect 511408 437376 511464 437410
rect 511498 437376 511554 437410
rect 511588 437376 511644 437410
rect 511678 437376 511734 437410
rect 511768 437376 511824 437410
rect 511858 437376 511914 437410
rect 511948 437376 512004 437410
rect 512038 437376 512094 437410
rect 512128 437376 512662 437410
rect 512696 437376 512752 437410
rect 512786 437376 512842 437410
rect 512876 437376 512932 437410
rect 512966 437376 513022 437410
rect 513056 437376 513112 437410
rect 513146 437376 513202 437410
rect 513236 437376 513292 437410
rect 513326 437376 513382 437410
rect 513416 437376 513674 437410
rect 503370 437362 513674 437376
rect 503370 437328 503402 437362
rect 503436 437328 504589 437362
rect 504623 437328 504690 437362
rect 504724 437328 505877 437362
rect 505911 437328 505978 437362
rect 506012 437328 507165 437362
rect 507199 437328 507266 437362
rect 507300 437328 508453 437362
rect 508487 437328 508554 437362
rect 508588 437328 509741 437362
rect 509775 437328 509842 437362
rect 509876 437328 511029 437362
rect 511063 437328 511130 437362
rect 511164 437328 512317 437362
rect 512351 437328 512418 437362
rect 512452 437328 513605 437362
rect 513639 437328 513674 437362
rect 503370 437261 513674 437328
rect 503370 437227 503486 437261
rect 503520 437227 503576 437261
rect 503610 437227 503666 437261
rect 503700 437227 503756 437261
rect 503790 437227 503846 437261
rect 503880 437227 503936 437261
rect 503970 437227 504026 437261
rect 504060 437227 504116 437261
rect 504150 437227 504206 437261
rect 504240 437227 504296 437261
rect 504330 437227 504386 437261
rect 504420 437227 504476 437261
rect 504510 437227 504566 437261
rect 504600 437227 504774 437261
rect 504808 437227 504864 437261
rect 504898 437227 504954 437261
rect 504988 437227 505044 437261
rect 505078 437227 505134 437261
rect 505168 437227 505224 437261
rect 505258 437227 505314 437261
rect 505348 437227 505404 437261
rect 505438 437227 505494 437261
rect 505528 437227 505584 437261
rect 505618 437227 505674 437261
rect 505708 437227 505764 437261
rect 505798 437227 505854 437261
rect 505888 437227 506062 437261
rect 506096 437227 506152 437261
rect 506186 437227 506242 437261
rect 506276 437227 506332 437261
rect 506366 437227 506422 437261
rect 506456 437227 506512 437261
rect 506546 437227 506602 437261
rect 506636 437227 506692 437261
rect 506726 437227 506782 437261
rect 506816 437227 506872 437261
rect 506906 437227 506962 437261
rect 506996 437227 507052 437261
rect 507086 437227 507142 437261
rect 507176 437227 507350 437261
rect 507384 437227 507440 437261
rect 507474 437227 507530 437261
rect 507564 437227 507620 437261
rect 507654 437227 507710 437261
rect 507744 437227 507800 437261
rect 507834 437227 507890 437261
rect 507924 437227 507980 437261
rect 508014 437227 508070 437261
rect 508104 437227 508160 437261
rect 508194 437227 508250 437261
rect 508284 437227 508340 437261
rect 508374 437227 508430 437261
rect 508464 437227 508638 437261
rect 508672 437227 508728 437261
rect 508762 437227 508818 437261
rect 508852 437227 508908 437261
rect 508942 437227 508998 437261
rect 509032 437227 509088 437261
rect 509122 437227 509178 437261
rect 509212 437227 509268 437261
rect 509302 437227 509358 437261
rect 509392 437227 509448 437261
rect 509482 437227 509538 437261
rect 509572 437227 509628 437261
rect 509662 437227 509718 437261
rect 509752 437227 509926 437261
rect 509960 437227 510016 437261
rect 510050 437227 510106 437261
rect 510140 437227 510196 437261
rect 510230 437227 510286 437261
rect 510320 437227 510376 437261
rect 510410 437227 510466 437261
rect 510500 437227 510556 437261
rect 510590 437227 510646 437261
rect 510680 437227 510736 437261
rect 510770 437227 510826 437261
rect 510860 437227 510916 437261
rect 510950 437227 511006 437261
rect 511040 437227 511214 437261
rect 511248 437227 511304 437261
rect 511338 437227 511394 437261
rect 511428 437227 511484 437261
rect 511518 437227 511574 437261
rect 511608 437227 511664 437261
rect 511698 437227 511754 437261
rect 511788 437227 511844 437261
rect 511878 437227 511934 437261
rect 511968 437227 512024 437261
rect 512058 437227 512114 437261
rect 512148 437227 512204 437261
rect 512238 437227 512294 437261
rect 512328 437227 512502 437261
rect 512536 437227 512592 437261
rect 512626 437227 512682 437261
rect 512716 437227 512772 437261
rect 512806 437227 512862 437261
rect 512896 437227 512952 437261
rect 512986 437227 513042 437261
rect 513076 437227 513132 437261
rect 513166 437227 513222 437261
rect 513256 437227 513312 437261
rect 513346 437227 513402 437261
rect 513436 437227 513492 437261
rect 513526 437227 513582 437261
rect 513616 437227 513674 437261
rect 501368 437092 501384 437216
rect 503370 437160 513674 437227
rect 516190 437832 516622 438046
rect 522926 437832 523358 438046
rect 516190 437816 523358 437832
rect 516190 437246 516622 437816
rect 522926 437246 523358 437816
rect 516190 437230 523358 437246
rect 516190 437222 516622 437230
rect 522926 437222 523358 437230
rect 503370 437126 503486 437160
rect 503520 437126 503576 437160
rect 503610 437126 503666 437160
rect 503700 437126 503756 437160
rect 503790 437126 503846 437160
rect 503880 437126 503936 437160
rect 503970 437126 504026 437160
rect 504060 437126 504116 437160
rect 504150 437126 504206 437160
rect 504240 437126 504296 437160
rect 504330 437126 504386 437160
rect 504420 437126 504476 437160
rect 504510 437126 504566 437160
rect 504600 437126 504774 437160
rect 504808 437126 504864 437160
rect 504898 437126 504954 437160
rect 504988 437126 505044 437160
rect 505078 437126 505134 437160
rect 505168 437126 505224 437160
rect 505258 437126 505314 437160
rect 505348 437126 505404 437160
rect 505438 437126 505494 437160
rect 505528 437126 505584 437160
rect 505618 437126 505674 437160
rect 505708 437126 505764 437160
rect 505798 437126 505854 437160
rect 505888 437126 506062 437160
rect 506096 437126 506152 437160
rect 506186 437126 506242 437160
rect 506276 437126 506332 437160
rect 506366 437126 506422 437160
rect 506456 437126 506512 437160
rect 506546 437126 506602 437160
rect 506636 437126 506692 437160
rect 506726 437126 506782 437160
rect 506816 437126 506872 437160
rect 506906 437126 506962 437160
rect 506996 437126 507052 437160
rect 507086 437126 507142 437160
rect 507176 437126 507350 437160
rect 507384 437126 507440 437160
rect 507474 437126 507530 437160
rect 507564 437126 507620 437160
rect 507654 437126 507710 437160
rect 507744 437126 507800 437160
rect 507834 437126 507890 437160
rect 507924 437126 507980 437160
rect 508014 437126 508070 437160
rect 508104 437126 508160 437160
rect 508194 437126 508250 437160
rect 508284 437126 508340 437160
rect 508374 437126 508430 437160
rect 508464 437126 508638 437160
rect 508672 437126 508728 437160
rect 508762 437126 508818 437160
rect 508852 437126 508908 437160
rect 508942 437126 508998 437160
rect 509032 437126 509088 437160
rect 509122 437126 509178 437160
rect 509212 437126 509268 437160
rect 509302 437126 509358 437160
rect 509392 437126 509448 437160
rect 509482 437126 509538 437160
rect 509572 437126 509628 437160
rect 509662 437126 509718 437160
rect 509752 437126 509926 437160
rect 509960 437126 510016 437160
rect 510050 437126 510106 437160
rect 510140 437126 510196 437160
rect 510230 437126 510286 437160
rect 510320 437126 510376 437160
rect 510410 437126 510466 437160
rect 510500 437126 510556 437160
rect 510590 437126 510646 437160
rect 510680 437126 510736 437160
rect 510770 437126 510826 437160
rect 510860 437126 510916 437160
rect 510950 437126 511006 437160
rect 511040 437126 511214 437160
rect 511248 437126 511304 437160
rect 511338 437126 511394 437160
rect 511428 437126 511484 437160
rect 511518 437126 511574 437160
rect 511608 437126 511664 437160
rect 511698 437126 511754 437160
rect 511788 437126 511844 437160
rect 511878 437126 511934 437160
rect 511968 437126 512024 437160
rect 512058 437126 512114 437160
rect 512148 437126 512204 437160
rect 512238 437126 512294 437160
rect 512328 437126 512502 437160
rect 512536 437126 512592 437160
rect 512626 437126 512682 437160
rect 512716 437126 512772 437160
rect 512806 437126 512862 437160
rect 512896 437126 512952 437160
rect 512986 437126 513042 437160
rect 513076 437126 513132 437160
rect 513166 437126 513222 437160
rect 513256 437126 513312 437160
rect 513346 437126 513402 437160
rect 513436 437126 513492 437160
rect 513526 437126 513582 437160
rect 513616 437126 513674 437160
rect 503370 437064 513674 437126
rect 503370 437030 503402 437064
rect 503436 437030 504589 437064
rect 504623 437030 504690 437064
rect 504724 437030 505877 437064
rect 505911 437030 505978 437064
rect 506012 437030 507165 437064
rect 507199 437030 507266 437064
rect 507300 437030 508453 437064
rect 508487 437030 508554 437064
rect 508588 437030 509741 437064
rect 509775 437030 509842 437064
rect 509876 437030 511029 437064
rect 511063 437030 511130 437064
rect 511164 437030 512317 437064
rect 512351 437030 512418 437064
rect 512452 437030 513605 437064
rect 513639 437030 513674 437064
rect 503370 437012 513674 437030
rect 501368 436868 501384 436992
rect 503370 436978 503665 437012
rect 503699 436978 503755 437012
rect 503789 436978 503845 437012
rect 503879 436978 503935 437012
rect 503969 436978 504025 437012
rect 504059 436978 504115 437012
rect 504149 436978 504205 437012
rect 504239 436978 504295 437012
rect 504329 436978 504385 437012
rect 504419 436978 504953 437012
rect 504987 436978 505043 437012
rect 505077 436978 505133 437012
rect 505167 436978 505223 437012
rect 505257 436978 505313 437012
rect 505347 436978 505403 437012
rect 505437 436978 505493 437012
rect 505527 436978 505583 437012
rect 505617 436978 505673 437012
rect 505707 436978 506241 437012
rect 506275 436978 506331 437012
rect 506365 436978 506421 437012
rect 506455 436978 506511 437012
rect 506545 436978 506601 437012
rect 506635 436978 506691 437012
rect 506725 436978 506781 437012
rect 506815 436978 506871 437012
rect 506905 436978 506961 437012
rect 506995 436978 507529 437012
rect 507563 436978 507619 437012
rect 507653 436978 507709 437012
rect 507743 436978 507799 437012
rect 507833 436978 507889 437012
rect 507923 436978 507979 437012
rect 508013 436978 508069 437012
rect 508103 436978 508159 437012
rect 508193 436978 508249 437012
rect 508283 436978 508817 437012
rect 508851 436978 508907 437012
rect 508941 436978 508997 437012
rect 509031 436978 509087 437012
rect 509121 436978 509177 437012
rect 509211 436978 509267 437012
rect 509301 436978 509357 437012
rect 509391 436978 509447 437012
rect 509481 436978 509537 437012
rect 509571 436978 510105 437012
rect 510139 436978 510195 437012
rect 510229 436978 510285 437012
rect 510319 436978 510375 437012
rect 510409 436978 510465 437012
rect 510499 436978 510555 437012
rect 510589 436978 510645 437012
rect 510679 436978 510735 437012
rect 510769 436978 510825 437012
rect 510859 436978 511393 437012
rect 511427 436978 511483 437012
rect 511517 436978 511573 437012
rect 511607 436978 511663 437012
rect 511697 436978 511753 437012
rect 511787 436978 511843 437012
rect 511877 436978 511933 437012
rect 511967 436978 512023 437012
rect 512057 436978 512113 437012
rect 512147 436978 512681 437012
rect 512715 436978 512771 437012
rect 512805 436978 512861 437012
rect 512895 436978 512951 437012
rect 512985 436978 513041 437012
rect 513075 436978 513131 437012
rect 513165 436978 513221 437012
rect 513255 436978 513311 437012
rect 513345 436978 513401 437012
rect 513435 436978 513674 437012
rect 503370 436974 513674 436978
rect 503370 436940 503402 436974
rect 503436 436959 504589 436974
rect 503436 436940 503605 436959
rect 503370 436934 503605 436940
rect 503370 436900 503552 436934
rect 503586 436900 503605 436934
rect 503370 436884 503605 436900
rect 504423 436940 504589 436959
rect 504623 436940 504690 436974
rect 504724 436959 505877 436974
rect 504724 436940 504893 436959
rect 504423 436934 504893 436940
rect 504423 436900 504840 436934
rect 504874 436900 504893 436934
rect 503370 436850 503402 436884
rect 503436 436850 503605 436884
rect 503370 436844 503605 436850
rect 503370 436810 503552 436844
rect 503586 436810 503605 436844
rect 503370 436794 503605 436810
rect 501368 436644 501384 436768
rect 503370 436760 503402 436794
rect 503436 436760 503605 436794
rect 503370 436754 503605 436760
rect 503370 436720 503552 436754
rect 503586 436720 503605 436754
rect 503370 436704 503605 436720
rect 503370 436670 503402 436704
rect 503436 436670 503605 436704
rect 503370 436664 503605 436670
rect 503370 436630 503552 436664
rect 503586 436630 503605 436664
rect 503370 436614 503605 436630
rect 503370 436580 503402 436614
rect 503436 436580 503605 436614
rect 503370 436574 503605 436580
rect 501368 436420 501384 436544
rect 503370 436540 503552 436574
rect 503586 436540 503605 436574
rect 503370 436524 503605 436540
rect 503370 436490 503402 436524
rect 503436 436490 503605 436524
rect 503370 436484 503605 436490
rect 503370 436450 503552 436484
rect 503586 436450 503605 436484
rect 503370 436434 503605 436450
rect 503370 436400 503402 436434
rect 503436 436400 503605 436434
rect 503370 436394 503605 436400
rect 503370 436360 503552 436394
rect 503586 436360 503605 436394
rect 503370 436344 503605 436360
rect 501368 436196 501384 436320
rect 503370 436310 503402 436344
rect 503436 436310 503605 436344
rect 503370 436304 503605 436310
rect 503370 436270 503552 436304
rect 503586 436270 503605 436304
rect 503370 436254 503605 436270
rect 503370 436220 503402 436254
rect 503436 436220 503605 436254
rect 503370 436214 503605 436220
rect 503370 436180 503552 436214
rect 503586 436180 503605 436214
rect 503667 436836 504361 436897
rect 503667 436802 503728 436836
rect 503762 436824 503818 436836
rect 503852 436824 503908 436836
rect 503942 436824 503998 436836
rect 503774 436802 503818 436824
rect 503874 436802 503908 436824
rect 503974 436802 503998 436824
rect 504032 436824 504088 436836
rect 504032 436802 504040 436824
rect 503667 436790 503740 436802
rect 503774 436790 503840 436802
rect 503874 436790 503940 436802
rect 503974 436790 504040 436802
rect 504074 436802 504088 436824
rect 504122 436824 504178 436836
rect 504122 436802 504140 436824
rect 504074 436790 504140 436802
rect 504174 436802 504178 436824
rect 504212 436824 504268 436836
rect 504212 436802 504240 436824
rect 504302 436802 504361 436836
rect 504174 436790 504240 436802
rect 504274 436790 504361 436802
rect 503667 436746 504361 436790
rect 503667 436712 503728 436746
rect 503762 436724 503818 436746
rect 503852 436724 503908 436746
rect 503942 436724 503998 436746
rect 503774 436712 503818 436724
rect 503874 436712 503908 436724
rect 503974 436712 503998 436724
rect 504032 436724 504088 436746
rect 504032 436712 504040 436724
rect 503667 436690 503740 436712
rect 503774 436690 503840 436712
rect 503874 436690 503940 436712
rect 503974 436690 504040 436712
rect 504074 436712 504088 436724
rect 504122 436724 504178 436746
rect 504122 436712 504140 436724
rect 504074 436690 504140 436712
rect 504174 436712 504178 436724
rect 504212 436724 504268 436746
rect 504212 436712 504240 436724
rect 504302 436712 504361 436746
rect 504174 436690 504240 436712
rect 504274 436690 504361 436712
rect 503667 436656 504361 436690
rect 503667 436622 503728 436656
rect 503762 436624 503818 436656
rect 503852 436624 503908 436656
rect 503942 436624 503998 436656
rect 503774 436622 503818 436624
rect 503874 436622 503908 436624
rect 503974 436622 503998 436624
rect 504032 436624 504088 436656
rect 504032 436622 504040 436624
rect 503667 436590 503740 436622
rect 503774 436590 503840 436622
rect 503874 436590 503940 436622
rect 503974 436590 504040 436622
rect 504074 436622 504088 436624
rect 504122 436624 504178 436656
rect 504122 436622 504140 436624
rect 504074 436590 504140 436622
rect 504174 436622 504178 436624
rect 504212 436624 504268 436656
rect 504212 436622 504240 436624
rect 504302 436622 504361 436656
rect 504174 436590 504240 436622
rect 504274 436590 504361 436622
rect 503667 436566 504361 436590
rect 503667 436532 503728 436566
rect 503762 436532 503818 436566
rect 503852 436532 503908 436566
rect 503942 436532 503998 436566
rect 504032 436532 504088 436566
rect 504122 436532 504178 436566
rect 504212 436532 504268 436566
rect 504302 436532 504361 436566
rect 503667 436524 504361 436532
rect 503667 436490 503740 436524
rect 503774 436490 503840 436524
rect 503874 436490 503940 436524
rect 503974 436490 504040 436524
rect 504074 436490 504140 436524
rect 504174 436490 504240 436524
rect 504274 436490 504361 436524
rect 503667 436476 504361 436490
rect 503667 436442 503728 436476
rect 503762 436442 503818 436476
rect 503852 436442 503908 436476
rect 503942 436442 503998 436476
rect 504032 436442 504088 436476
rect 504122 436442 504178 436476
rect 504212 436442 504268 436476
rect 504302 436442 504361 436476
rect 503667 436424 504361 436442
rect 503667 436390 503740 436424
rect 503774 436390 503840 436424
rect 503874 436390 503940 436424
rect 503974 436390 504040 436424
rect 504074 436390 504140 436424
rect 504174 436390 504240 436424
rect 504274 436390 504361 436424
rect 503667 436386 504361 436390
rect 503667 436352 503728 436386
rect 503762 436352 503818 436386
rect 503852 436352 503908 436386
rect 503942 436352 503998 436386
rect 504032 436352 504088 436386
rect 504122 436352 504178 436386
rect 504212 436352 504268 436386
rect 504302 436352 504361 436386
rect 503667 436324 504361 436352
rect 503667 436296 503740 436324
rect 503774 436296 503840 436324
rect 503874 436296 503940 436324
rect 503974 436296 504040 436324
rect 503667 436262 503728 436296
rect 503774 436290 503818 436296
rect 503874 436290 503908 436296
rect 503974 436290 503998 436296
rect 503762 436262 503818 436290
rect 503852 436262 503908 436290
rect 503942 436262 503998 436290
rect 504032 436290 504040 436296
rect 504074 436296 504140 436324
rect 504074 436290 504088 436296
rect 504032 436262 504088 436290
rect 504122 436290 504140 436296
rect 504174 436296 504240 436324
rect 504274 436296 504361 436324
rect 504174 436290 504178 436296
rect 504122 436262 504178 436290
rect 504212 436290 504240 436296
rect 504212 436262 504268 436290
rect 504302 436262 504361 436296
rect 503667 436203 504361 436262
rect 504423 436866 504442 436900
rect 504476 436884 504893 436900
rect 505711 436940 505877 436959
rect 505911 436940 505978 436974
rect 506012 436959 507165 436974
rect 506012 436940 506181 436959
rect 505711 436934 506181 436940
rect 505711 436900 506128 436934
rect 506162 436900 506181 436934
rect 504476 436866 504589 436884
rect 504423 436850 504589 436866
rect 504623 436850 504690 436884
rect 504724 436850 504893 436884
rect 504423 436844 504893 436850
rect 504423 436810 504840 436844
rect 504874 436810 504893 436844
rect 504423 436776 504442 436810
rect 504476 436794 504893 436810
rect 504476 436776 504589 436794
rect 504423 436760 504589 436776
rect 504623 436760 504690 436794
rect 504724 436760 504893 436794
rect 504423 436754 504893 436760
rect 504423 436720 504840 436754
rect 504874 436720 504893 436754
rect 504423 436686 504442 436720
rect 504476 436704 504893 436720
rect 504476 436686 504589 436704
rect 504423 436670 504589 436686
rect 504623 436670 504690 436704
rect 504724 436670 504893 436704
rect 504423 436664 504893 436670
rect 504423 436630 504840 436664
rect 504874 436630 504893 436664
rect 504423 436596 504442 436630
rect 504476 436614 504893 436630
rect 504476 436596 504589 436614
rect 504423 436580 504589 436596
rect 504623 436580 504690 436614
rect 504724 436580 504893 436614
rect 504423 436574 504893 436580
rect 504423 436540 504840 436574
rect 504874 436540 504893 436574
rect 504423 436506 504442 436540
rect 504476 436524 504893 436540
rect 504476 436506 504589 436524
rect 504423 436490 504589 436506
rect 504623 436490 504690 436524
rect 504724 436490 504893 436524
rect 504423 436484 504893 436490
rect 504423 436450 504840 436484
rect 504874 436450 504893 436484
rect 504423 436416 504442 436450
rect 504476 436434 504893 436450
rect 504476 436416 504589 436434
rect 504423 436400 504589 436416
rect 504623 436400 504690 436434
rect 504724 436400 504893 436434
rect 504423 436394 504893 436400
rect 504423 436360 504840 436394
rect 504874 436360 504893 436394
rect 504423 436326 504442 436360
rect 504476 436344 504893 436360
rect 504476 436326 504589 436344
rect 504423 436310 504589 436326
rect 504623 436310 504690 436344
rect 504724 436310 504893 436344
rect 504423 436304 504893 436310
rect 504423 436270 504840 436304
rect 504874 436270 504893 436304
rect 504423 436236 504442 436270
rect 504476 436254 504893 436270
rect 504476 436236 504589 436254
rect 504423 436220 504589 436236
rect 504623 436220 504690 436254
rect 504724 436220 504893 436254
rect 504423 436214 504893 436220
rect 503370 436164 503605 436180
rect 503370 436130 503402 436164
rect 503436 436141 503605 436164
rect 504423 436180 504840 436214
rect 504874 436180 504893 436214
rect 504955 436836 505649 436897
rect 504955 436802 505016 436836
rect 505050 436824 505106 436836
rect 505140 436824 505196 436836
rect 505230 436824 505286 436836
rect 505062 436802 505106 436824
rect 505162 436802 505196 436824
rect 505262 436802 505286 436824
rect 505320 436824 505376 436836
rect 505320 436802 505328 436824
rect 504955 436790 505028 436802
rect 505062 436790 505128 436802
rect 505162 436790 505228 436802
rect 505262 436790 505328 436802
rect 505362 436802 505376 436824
rect 505410 436824 505466 436836
rect 505410 436802 505428 436824
rect 505362 436790 505428 436802
rect 505462 436802 505466 436824
rect 505500 436824 505556 436836
rect 505500 436802 505528 436824
rect 505590 436802 505649 436836
rect 505462 436790 505528 436802
rect 505562 436790 505649 436802
rect 504955 436746 505649 436790
rect 504955 436712 505016 436746
rect 505050 436724 505106 436746
rect 505140 436724 505196 436746
rect 505230 436724 505286 436746
rect 505062 436712 505106 436724
rect 505162 436712 505196 436724
rect 505262 436712 505286 436724
rect 505320 436724 505376 436746
rect 505320 436712 505328 436724
rect 504955 436690 505028 436712
rect 505062 436690 505128 436712
rect 505162 436690 505228 436712
rect 505262 436690 505328 436712
rect 505362 436712 505376 436724
rect 505410 436724 505466 436746
rect 505410 436712 505428 436724
rect 505362 436690 505428 436712
rect 505462 436712 505466 436724
rect 505500 436724 505556 436746
rect 505500 436712 505528 436724
rect 505590 436712 505649 436746
rect 505462 436690 505528 436712
rect 505562 436690 505649 436712
rect 504955 436656 505649 436690
rect 504955 436622 505016 436656
rect 505050 436624 505106 436656
rect 505140 436624 505196 436656
rect 505230 436624 505286 436656
rect 505062 436622 505106 436624
rect 505162 436622 505196 436624
rect 505262 436622 505286 436624
rect 505320 436624 505376 436656
rect 505320 436622 505328 436624
rect 504955 436590 505028 436622
rect 505062 436590 505128 436622
rect 505162 436590 505228 436622
rect 505262 436590 505328 436622
rect 505362 436622 505376 436624
rect 505410 436624 505466 436656
rect 505410 436622 505428 436624
rect 505362 436590 505428 436622
rect 505462 436622 505466 436624
rect 505500 436624 505556 436656
rect 505500 436622 505528 436624
rect 505590 436622 505649 436656
rect 505462 436590 505528 436622
rect 505562 436590 505649 436622
rect 504955 436566 505649 436590
rect 504955 436532 505016 436566
rect 505050 436532 505106 436566
rect 505140 436532 505196 436566
rect 505230 436532 505286 436566
rect 505320 436532 505376 436566
rect 505410 436532 505466 436566
rect 505500 436532 505556 436566
rect 505590 436532 505649 436566
rect 504955 436524 505649 436532
rect 504955 436490 505028 436524
rect 505062 436490 505128 436524
rect 505162 436490 505228 436524
rect 505262 436490 505328 436524
rect 505362 436490 505428 436524
rect 505462 436490 505528 436524
rect 505562 436490 505649 436524
rect 504955 436476 505649 436490
rect 504955 436442 505016 436476
rect 505050 436442 505106 436476
rect 505140 436442 505196 436476
rect 505230 436442 505286 436476
rect 505320 436442 505376 436476
rect 505410 436442 505466 436476
rect 505500 436442 505556 436476
rect 505590 436442 505649 436476
rect 504955 436424 505649 436442
rect 504955 436390 505028 436424
rect 505062 436390 505128 436424
rect 505162 436390 505228 436424
rect 505262 436390 505328 436424
rect 505362 436390 505428 436424
rect 505462 436390 505528 436424
rect 505562 436390 505649 436424
rect 504955 436386 505649 436390
rect 504955 436352 505016 436386
rect 505050 436352 505106 436386
rect 505140 436352 505196 436386
rect 505230 436352 505286 436386
rect 505320 436352 505376 436386
rect 505410 436352 505466 436386
rect 505500 436352 505556 436386
rect 505590 436352 505649 436386
rect 504955 436324 505649 436352
rect 504955 436296 505028 436324
rect 505062 436296 505128 436324
rect 505162 436296 505228 436324
rect 505262 436296 505328 436324
rect 504955 436262 505016 436296
rect 505062 436290 505106 436296
rect 505162 436290 505196 436296
rect 505262 436290 505286 436296
rect 505050 436262 505106 436290
rect 505140 436262 505196 436290
rect 505230 436262 505286 436290
rect 505320 436290 505328 436296
rect 505362 436296 505428 436324
rect 505362 436290 505376 436296
rect 505320 436262 505376 436290
rect 505410 436290 505428 436296
rect 505462 436296 505528 436324
rect 505562 436296 505649 436324
rect 505462 436290 505466 436296
rect 505410 436262 505466 436290
rect 505500 436290 505528 436296
rect 505500 436262 505556 436290
rect 505590 436262 505649 436296
rect 504955 436203 505649 436262
rect 505711 436866 505730 436900
rect 505764 436884 506181 436900
rect 506999 436940 507165 436959
rect 507199 436940 507266 436974
rect 507300 436959 508453 436974
rect 507300 436940 507469 436959
rect 506999 436934 507469 436940
rect 506999 436900 507416 436934
rect 507450 436900 507469 436934
rect 505764 436866 505877 436884
rect 505711 436850 505877 436866
rect 505911 436850 505978 436884
rect 506012 436850 506181 436884
rect 505711 436844 506181 436850
rect 505711 436810 506128 436844
rect 506162 436810 506181 436844
rect 505711 436776 505730 436810
rect 505764 436794 506181 436810
rect 505764 436776 505877 436794
rect 505711 436760 505877 436776
rect 505911 436760 505978 436794
rect 506012 436760 506181 436794
rect 505711 436754 506181 436760
rect 505711 436720 506128 436754
rect 506162 436720 506181 436754
rect 505711 436686 505730 436720
rect 505764 436704 506181 436720
rect 505764 436686 505877 436704
rect 505711 436670 505877 436686
rect 505911 436670 505978 436704
rect 506012 436670 506181 436704
rect 505711 436664 506181 436670
rect 505711 436630 506128 436664
rect 506162 436630 506181 436664
rect 505711 436596 505730 436630
rect 505764 436614 506181 436630
rect 505764 436596 505877 436614
rect 505711 436580 505877 436596
rect 505911 436580 505978 436614
rect 506012 436580 506181 436614
rect 505711 436574 506181 436580
rect 505711 436540 506128 436574
rect 506162 436540 506181 436574
rect 505711 436506 505730 436540
rect 505764 436524 506181 436540
rect 505764 436506 505877 436524
rect 505711 436490 505877 436506
rect 505911 436490 505978 436524
rect 506012 436490 506181 436524
rect 505711 436484 506181 436490
rect 505711 436450 506128 436484
rect 506162 436450 506181 436484
rect 505711 436416 505730 436450
rect 505764 436434 506181 436450
rect 505764 436416 505877 436434
rect 505711 436400 505877 436416
rect 505911 436400 505978 436434
rect 506012 436400 506181 436434
rect 505711 436394 506181 436400
rect 505711 436360 506128 436394
rect 506162 436360 506181 436394
rect 505711 436326 505730 436360
rect 505764 436344 506181 436360
rect 505764 436326 505877 436344
rect 505711 436310 505877 436326
rect 505911 436310 505978 436344
rect 506012 436310 506181 436344
rect 505711 436304 506181 436310
rect 505711 436270 506128 436304
rect 506162 436270 506181 436304
rect 505711 436236 505730 436270
rect 505764 436254 506181 436270
rect 505764 436236 505877 436254
rect 505711 436220 505877 436236
rect 505911 436220 505978 436254
rect 506012 436220 506181 436254
rect 505711 436214 506181 436220
rect 504423 436146 504442 436180
rect 504476 436164 504893 436180
rect 504476 436146 504589 436164
rect 504423 436141 504589 436146
rect 503436 436130 504589 436141
rect 504623 436130 504690 436164
rect 504724 436141 504893 436164
rect 505711 436180 506128 436214
rect 506162 436180 506181 436214
rect 506243 436836 506937 436897
rect 506243 436802 506304 436836
rect 506338 436824 506394 436836
rect 506428 436824 506484 436836
rect 506518 436824 506574 436836
rect 506350 436802 506394 436824
rect 506450 436802 506484 436824
rect 506550 436802 506574 436824
rect 506608 436824 506664 436836
rect 506608 436802 506616 436824
rect 506243 436790 506316 436802
rect 506350 436790 506416 436802
rect 506450 436790 506516 436802
rect 506550 436790 506616 436802
rect 506650 436802 506664 436824
rect 506698 436824 506754 436836
rect 506698 436802 506716 436824
rect 506650 436790 506716 436802
rect 506750 436802 506754 436824
rect 506788 436824 506844 436836
rect 506788 436802 506816 436824
rect 506878 436802 506937 436836
rect 506750 436790 506816 436802
rect 506850 436790 506937 436802
rect 506243 436746 506937 436790
rect 506243 436712 506304 436746
rect 506338 436724 506394 436746
rect 506428 436724 506484 436746
rect 506518 436724 506574 436746
rect 506350 436712 506394 436724
rect 506450 436712 506484 436724
rect 506550 436712 506574 436724
rect 506608 436724 506664 436746
rect 506608 436712 506616 436724
rect 506243 436690 506316 436712
rect 506350 436690 506416 436712
rect 506450 436690 506516 436712
rect 506550 436690 506616 436712
rect 506650 436712 506664 436724
rect 506698 436724 506754 436746
rect 506698 436712 506716 436724
rect 506650 436690 506716 436712
rect 506750 436712 506754 436724
rect 506788 436724 506844 436746
rect 506788 436712 506816 436724
rect 506878 436712 506937 436746
rect 506750 436690 506816 436712
rect 506850 436690 506937 436712
rect 506243 436656 506937 436690
rect 506243 436622 506304 436656
rect 506338 436624 506394 436656
rect 506428 436624 506484 436656
rect 506518 436624 506574 436656
rect 506350 436622 506394 436624
rect 506450 436622 506484 436624
rect 506550 436622 506574 436624
rect 506608 436624 506664 436656
rect 506608 436622 506616 436624
rect 506243 436590 506316 436622
rect 506350 436590 506416 436622
rect 506450 436590 506516 436622
rect 506550 436590 506616 436622
rect 506650 436622 506664 436624
rect 506698 436624 506754 436656
rect 506698 436622 506716 436624
rect 506650 436590 506716 436622
rect 506750 436622 506754 436624
rect 506788 436624 506844 436656
rect 506788 436622 506816 436624
rect 506878 436622 506937 436656
rect 506750 436590 506816 436622
rect 506850 436590 506937 436622
rect 506243 436566 506937 436590
rect 506243 436532 506304 436566
rect 506338 436532 506394 436566
rect 506428 436532 506484 436566
rect 506518 436532 506574 436566
rect 506608 436532 506664 436566
rect 506698 436532 506754 436566
rect 506788 436532 506844 436566
rect 506878 436532 506937 436566
rect 506243 436524 506937 436532
rect 506243 436490 506316 436524
rect 506350 436490 506416 436524
rect 506450 436490 506516 436524
rect 506550 436490 506616 436524
rect 506650 436490 506716 436524
rect 506750 436490 506816 436524
rect 506850 436490 506937 436524
rect 506243 436476 506937 436490
rect 506243 436442 506304 436476
rect 506338 436442 506394 436476
rect 506428 436442 506484 436476
rect 506518 436442 506574 436476
rect 506608 436442 506664 436476
rect 506698 436442 506754 436476
rect 506788 436442 506844 436476
rect 506878 436442 506937 436476
rect 506243 436424 506937 436442
rect 506243 436390 506316 436424
rect 506350 436390 506416 436424
rect 506450 436390 506516 436424
rect 506550 436390 506616 436424
rect 506650 436390 506716 436424
rect 506750 436390 506816 436424
rect 506850 436390 506937 436424
rect 506243 436386 506937 436390
rect 506243 436352 506304 436386
rect 506338 436352 506394 436386
rect 506428 436352 506484 436386
rect 506518 436352 506574 436386
rect 506608 436352 506664 436386
rect 506698 436352 506754 436386
rect 506788 436352 506844 436386
rect 506878 436352 506937 436386
rect 506243 436324 506937 436352
rect 506243 436296 506316 436324
rect 506350 436296 506416 436324
rect 506450 436296 506516 436324
rect 506550 436296 506616 436324
rect 506243 436262 506304 436296
rect 506350 436290 506394 436296
rect 506450 436290 506484 436296
rect 506550 436290 506574 436296
rect 506338 436262 506394 436290
rect 506428 436262 506484 436290
rect 506518 436262 506574 436290
rect 506608 436290 506616 436296
rect 506650 436296 506716 436324
rect 506650 436290 506664 436296
rect 506608 436262 506664 436290
rect 506698 436290 506716 436296
rect 506750 436296 506816 436324
rect 506850 436296 506937 436324
rect 506750 436290 506754 436296
rect 506698 436262 506754 436290
rect 506788 436290 506816 436296
rect 506788 436262 506844 436290
rect 506878 436262 506937 436296
rect 506243 436203 506937 436262
rect 506999 436866 507018 436900
rect 507052 436884 507469 436900
rect 508287 436940 508453 436959
rect 508487 436940 508554 436974
rect 508588 436959 509741 436974
rect 508588 436940 508757 436959
rect 508287 436934 508757 436940
rect 508287 436900 508704 436934
rect 508738 436900 508757 436934
rect 507052 436866 507165 436884
rect 506999 436850 507165 436866
rect 507199 436850 507266 436884
rect 507300 436850 507469 436884
rect 506999 436844 507469 436850
rect 506999 436810 507416 436844
rect 507450 436810 507469 436844
rect 506999 436776 507018 436810
rect 507052 436794 507469 436810
rect 507052 436776 507165 436794
rect 506999 436760 507165 436776
rect 507199 436760 507266 436794
rect 507300 436760 507469 436794
rect 506999 436754 507469 436760
rect 506999 436720 507416 436754
rect 507450 436720 507469 436754
rect 506999 436686 507018 436720
rect 507052 436704 507469 436720
rect 507052 436686 507165 436704
rect 506999 436670 507165 436686
rect 507199 436670 507266 436704
rect 507300 436670 507469 436704
rect 506999 436664 507469 436670
rect 506999 436630 507416 436664
rect 507450 436630 507469 436664
rect 506999 436596 507018 436630
rect 507052 436614 507469 436630
rect 507052 436596 507165 436614
rect 506999 436580 507165 436596
rect 507199 436580 507266 436614
rect 507300 436580 507469 436614
rect 506999 436574 507469 436580
rect 506999 436540 507416 436574
rect 507450 436540 507469 436574
rect 506999 436506 507018 436540
rect 507052 436524 507469 436540
rect 507052 436506 507165 436524
rect 506999 436490 507165 436506
rect 507199 436490 507266 436524
rect 507300 436490 507469 436524
rect 506999 436484 507469 436490
rect 506999 436450 507416 436484
rect 507450 436450 507469 436484
rect 506999 436416 507018 436450
rect 507052 436434 507469 436450
rect 507052 436416 507165 436434
rect 506999 436400 507165 436416
rect 507199 436400 507266 436434
rect 507300 436400 507469 436434
rect 506999 436394 507469 436400
rect 506999 436360 507416 436394
rect 507450 436360 507469 436394
rect 506999 436326 507018 436360
rect 507052 436344 507469 436360
rect 507052 436326 507165 436344
rect 506999 436310 507165 436326
rect 507199 436310 507266 436344
rect 507300 436310 507469 436344
rect 506999 436304 507469 436310
rect 506999 436270 507416 436304
rect 507450 436270 507469 436304
rect 506999 436236 507018 436270
rect 507052 436254 507469 436270
rect 507052 436236 507165 436254
rect 506999 436220 507165 436236
rect 507199 436220 507266 436254
rect 507300 436220 507469 436254
rect 506999 436214 507469 436220
rect 505711 436146 505730 436180
rect 505764 436164 506181 436180
rect 505764 436146 505877 436164
rect 505711 436141 505877 436146
rect 504724 436130 505877 436141
rect 505911 436130 505978 436164
rect 506012 436141 506181 436164
rect 506999 436180 507416 436214
rect 507450 436180 507469 436214
rect 507531 436836 508225 436897
rect 507531 436802 507592 436836
rect 507626 436824 507682 436836
rect 507716 436824 507772 436836
rect 507806 436824 507862 436836
rect 507638 436802 507682 436824
rect 507738 436802 507772 436824
rect 507838 436802 507862 436824
rect 507896 436824 507952 436836
rect 507896 436802 507904 436824
rect 507531 436790 507604 436802
rect 507638 436790 507704 436802
rect 507738 436790 507804 436802
rect 507838 436790 507904 436802
rect 507938 436802 507952 436824
rect 507986 436824 508042 436836
rect 507986 436802 508004 436824
rect 507938 436790 508004 436802
rect 508038 436802 508042 436824
rect 508076 436824 508132 436836
rect 508076 436802 508104 436824
rect 508166 436802 508225 436836
rect 508038 436790 508104 436802
rect 508138 436790 508225 436802
rect 507531 436746 508225 436790
rect 507531 436712 507592 436746
rect 507626 436724 507682 436746
rect 507716 436724 507772 436746
rect 507806 436724 507862 436746
rect 507638 436712 507682 436724
rect 507738 436712 507772 436724
rect 507838 436712 507862 436724
rect 507896 436724 507952 436746
rect 507896 436712 507904 436724
rect 507531 436690 507604 436712
rect 507638 436690 507704 436712
rect 507738 436690 507804 436712
rect 507838 436690 507904 436712
rect 507938 436712 507952 436724
rect 507986 436724 508042 436746
rect 507986 436712 508004 436724
rect 507938 436690 508004 436712
rect 508038 436712 508042 436724
rect 508076 436724 508132 436746
rect 508076 436712 508104 436724
rect 508166 436712 508225 436746
rect 508038 436690 508104 436712
rect 508138 436690 508225 436712
rect 507531 436656 508225 436690
rect 507531 436622 507592 436656
rect 507626 436624 507682 436656
rect 507716 436624 507772 436656
rect 507806 436624 507862 436656
rect 507638 436622 507682 436624
rect 507738 436622 507772 436624
rect 507838 436622 507862 436624
rect 507896 436624 507952 436656
rect 507896 436622 507904 436624
rect 507531 436590 507604 436622
rect 507638 436590 507704 436622
rect 507738 436590 507804 436622
rect 507838 436590 507904 436622
rect 507938 436622 507952 436624
rect 507986 436624 508042 436656
rect 507986 436622 508004 436624
rect 507938 436590 508004 436622
rect 508038 436622 508042 436624
rect 508076 436624 508132 436656
rect 508076 436622 508104 436624
rect 508166 436622 508225 436656
rect 508038 436590 508104 436622
rect 508138 436590 508225 436622
rect 507531 436566 508225 436590
rect 507531 436532 507592 436566
rect 507626 436532 507682 436566
rect 507716 436532 507772 436566
rect 507806 436532 507862 436566
rect 507896 436532 507952 436566
rect 507986 436532 508042 436566
rect 508076 436532 508132 436566
rect 508166 436532 508225 436566
rect 507531 436524 508225 436532
rect 507531 436490 507604 436524
rect 507638 436490 507704 436524
rect 507738 436490 507804 436524
rect 507838 436490 507904 436524
rect 507938 436490 508004 436524
rect 508038 436490 508104 436524
rect 508138 436490 508225 436524
rect 507531 436476 508225 436490
rect 507531 436442 507592 436476
rect 507626 436442 507682 436476
rect 507716 436442 507772 436476
rect 507806 436442 507862 436476
rect 507896 436442 507952 436476
rect 507986 436442 508042 436476
rect 508076 436442 508132 436476
rect 508166 436442 508225 436476
rect 507531 436424 508225 436442
rect 507531 436390 507604 436424
rect 507638 436390 507704 436424
rect 507738 436390 507804 436424
rect 507838 436390 507904 436424
rect 507938 436390 508004 436424
rect 508038 436390 508104 436424
rect 508138 436390 508225 436424
rect 507531 436386 508225 436390
rect 507531 436352 507592 436386
rect 507626 436352 507682 436386
rect 507716 436352 507772 436386
rect 507806 436352 507862 436386
rect 507896 436352 507952 436386
rect 507986 436352 508042 436386
rect 508076 436352 508132 436386
rect 508166 436352 508225 436386
rect 507531 436324 508225 436352
rect 507531 436296 507604 436324
rect 507638 436296 507704 436324
rect 507738 436296 507804 436324
rect 507838 436296 507904 436324
rect 507531 436262 507592 436296
rect 507638 436290 507682 436296
rect 507738 436290 507772 436296
rect 507838 436290 507862 436296
rect 507626 436262 507682 436290
rect 507716 436262 507772 436290
rect 507806 436262 507862 436290
rect 507896 436290 507904 436296
rect 507938 436296 508004 436324
rect 507938 436290 507952 436296
rect 507896 436262 507952 436290
rect 507986 436290 508004 436296
rect 508038 436296 508104 436324
rect 508138 436296 508225 436324
rect 508038 436290 508042 436296
rect 507986 436262 508042 436290
rect 508076 436290 508104 436296
rect 508076 436262 508132 436290
rect 508166 436262 508225 436296
rect 507531 436203 508225 436262
rect 508287 436866 508306 436900
rect 508340 436884 508757 436900
rect 509575 436940 509741 436959
rect 509775 436940 509842 436974
rect 509876 436959 511029 436974
rect 509876 436940 510045 436959
rect 509575 436934 510045 436940
rect 509575 436900 509992 436934
rect 510026 436900 510045 436934
rect 508340 436866 508453 436884
rect 508287 436850 508453 436866
rect 508487 436850 508554 436884
rect 508588 436850 508757 436884
rect 508287 436844 508757 436850
rect 508287 436810 508704 436844
rect 508738 436810 508757 436844
rect 508287 436776 508306 436810
rect 508340 436794 508757 436810
rect 508340 436776 508453 436794
rect 508287 436760 508453 436776
rect 508487 436760 508554 436794
rect 508588 436760 508757 436794
rect 508287 436754 508757 436760
rect 508287 436720 508704 436754
rect 508738 436720 508757 436754
rect 508287 436686 508306 436720
rect 508340 436704 508757 436720
rect 508340 436686 508453 436704
rect 508287 436670 508453 436686
rect 508487 436670 508554 436704
rect 508588 436670 508757 436704
rect 508287 436664 508757 436670
rect 508287 436630 508704 436664
rect 508738 436630 508757 436664
rect 508287 436596 508306 436630
rect 508340 436614 508757 436630
rect 508340 436596 508453 436614
rect 508287 436580 508453 436596
rect 508487 436580 508554 436614
rect 508588 436580 508757 436614
rect 508287 436574 508757 436580
rect 508287 436540 508704 436574
rect 508738 436540 508757 436574
rect 508287 436506 508306 436540
rect 508340 436524 508757 436540
rect 508340 436506 508453 436524
rect 508287 436490 508453 436506
rect 508487 436490 508554 436524
rect 508588 436490 508757 436524
rect 508287 436484 508757 436490
rect 508287 436450 508704 436484
rect 508738 436450 508757 436484
rect 508287 436416 508306 436450
rect 508340 436434 508757 436450
rect 508340 436416 508453 436434
rect 508287 436400 508453 436416
rect 508487 436400 508554 436434
rect 508588 436400 508757 436434
rect 508287 436394 508757 436400
rect 508287 436360 508704 436394
rect 508738 436360 508757 436394
rect 508287 436326 508306 436360
rect 508340 436344 508757 436360
rect 508340 436326 508453 436344
rect 508287 436310 508453 436326
rect 508487 436310 508554 436344
rect 508588 436310 508757 436344
rect 508287 436304 508757 436310
rect 508287 436270 508704 436304
rect 508738 436270 508757 436304
rect 508287 436236 508306 436270
rect 508340 436254 508757 436270
rect 508340 436236 508453 436254
rect 508287 436220 508453 436236
rect 508487 436220 508554 436254
rect 508588 436220 508757 436254
rect 508287 436214 508757 436220
rect 506999 436146 507018 436180
rect 507052 436164 507469 436180
rect 507052 436146 507165 436164
rect 506999 436141 507165 436146
rect 506012 436130 507165 436141
rect 507199 436130 507266 436164
rect 507300 436141 507469 436164
rect 508287 436180 508704 436214
rect 508738 436180 508757 436214
rect 508819 436836 509513 436897
rect 508819 436802 508880 436836
rect 508914 436824 508970 436836
rect 509004 436824 509060 436836
rect 509094 436824 509150 436836
rect 508926 436802 508970 436824
rect 509026 436802 509060 436824
rect 509126 436802 509150 436824
rect 509184 436824 509240 436836
rect 509184 436802 509192 436824
rect 508819 436790 508892 436802
rect 508926 436790 508992 436802
rect 509026 436790 509092 436802
rect 509126 436790 509192 436802
rect 509226 436802 509240 436824
rect 509274 436824 509330 436836
rect 509274 436802 509292 436824
rect 509226 436790 509292 436802
rect 509326 436802 509330 436824
rect 509364 436824 509420 436836
rect 509364 436802 509392 436824
rect 509454 436802 509513 436836
rect 509326 436790 509392 436802
rect 509426 436790 509513 436802
rect 508819 436746 509513 436790
rect 508819 436712 508880 436746
rect 508914 436724 508970 436746
rect 509004 436724 509060 436746
rect 509094 436724 509150 436746
rect 508926 436712 508970 436724
rect 509026 436712 509060 436724
rect 509126 436712 509150 436724
rect 509184 436724 509240 436746
rect 509184 436712 509192 436724
rect 508819 436690 508892 436712
rect 508926 436690 508992 436712
rect 509026 436690 509092 436712
rect 509126 436690 509192 436712
rect 509226 436712 509240 436724
rect 509274 436724 509330 436746
rect 509274 436712 509292 436724
rect 509226 436690 509292 436712
rect 509326 436712 509330 436724
rect 509364 436724 509420 436746
rect 509364 436712 509392 436724
rect 509454 436712 509513 436746
rect 509326 436690 509392 436712
rect 509426 436690 509513 436712
rect 508819 436656 509513 436690
rect 508819 436622 508880 436656
rect 508914 436624 508970 436656
rect 509004 436624 509060 436656
rect 509094 436624 509150 436656
rect 508926 436622 508970 436624
rect 509026 436622 509060 436624
rect 509126 436622 509150 436624
rect 509184 436624 509240 436656
rect 509184 436622 509192 436624
rect 508819 436590 508892 436622
rect 508926 436590 508992 436622
rect 509026 436590 509092 436622
rect 509126 436590 509192 436622
rect 509226 436622 509240 436624
rect 509274 436624 509330 436656
rect 509274 436622 509292 436624
rect 509226 436590 509292 436622
rect 509326 436622 509330 436624
rect 509364 436624 509420 436656
rect 509364 436622 509392 436624
rect 509454 436622 509513 436656
rect 509326 436590 509392 436622
rect 509426 436590 509513 436622
rect 508819 436566 509513 436590
rect 508819 436532 508880 436566
rect 508914 436532 508970 436566
rect 509004 436532 509060 436566
rect 509094 436532 509150 436566
rect 509184 436532 509240 436566
rect 509274 436532 509330 436566
rect 509364 436532 509420 436566
rect 509454 436532 509513 436566
rect 508819 436524 509513 436532
rect 508819 436490 508892 436524
rect 508926 436490 508992 436524
rect 509026 436490 509092 436524
rect 509126 436490 509192 436524
rect 509226 436490 509292 436524
rect 509326 436490 509392 436524
rect 509426 436490 509513 436524
rect 508819 436476 509513 436490
rect 508819 436442 508880 436476
rect 508914 436442 508970 436476
rect 509004 436442 509060 436476
rect 509094 436442 509150 436476
rect 509184 436442 509240 436476
rect 509274 436442 509330 436476
rect 509364 436442 509420 436476
rect 509454 436442 509513 436476
rect 508819 436424 509513 436442
rect 508819 436390 508892 436424
rect 508926 436390 508992 436424
rect 509026 436390 509092 436424
rect 509126 436390 509192 436424
rect 509226 436390 509292 436424
rect 509326 436390 509392 436424
rect 509426 436390 509513 436424
rect 508819 436386 509513 436390
rect 508819 436352 508880 436386
rect 508914 436352 508970 436386
rect 509004 436352 509060 436386
rect 509094 436352 509150 436386
rect 509184 436352 509240 436386
rect 509274 436352 509330 436386
rect 509364 436352 509420 436386
rect 509454 436352 509513 436386
rect 508819 436324 509513 436352
rect 508819 436296 508892 436324
rect 508926 436296 508992 436324
rect 509026 436296 509092 436324
rect 509126 436296 509192 436324
rect 508819 436262 508880 436296
rect 508926 436290 508970 436296
rect 509026 436290 509060 436296
rect 509126 436290 509150 436296
rect 508914 436262 508970 436290
rect 509004 436262 509060 436290
rect 509094 436262 509150 436290
rect 509184 436290 509192 436296
rect 509226 436296 509292 436324
rect 509226 436290 509240 436296
rect 509184 436262 509240 436290
rect 509274 436290 509292 436296
rect 509326 436296 509392 436324
rect 509426 436296 509513 436324
rect 509326 436290 509330 436296
rect 509274 436262 509330 436290
rect 509364 436290 509392 436296
rect 509364 436262 509420 436290
rect 509454 436262 509513 436296
rect 508819 436203 509513 436262
rect 509575 436866 509594 436900
rect 509628 436884 510045 436900
rect 510863 436940 511029 436959
rect 511063 436940 511130 436974
rect 511164 436959 512317 436974
rect 511164 436940 511333 436959
rect 510863 436934 511333 436940
rect 510863 436900 511280 436934
rect 511314 436900 511333 436934
rect 509628 436866 509741 436884
rect 509575 436850 509741 436866
rect 509775 436850 509842 436884
rect 509876 436850 510045 436884
rect 509575 436844 510045 436850
rect 509575 436810 509992 436844
rect 510026 436810 510045 436844
rect 509575 436776 509594 436810
rect 509628 436794 510045 436810
rect 509628 436776 509741 436794
rect 509575 436760 509741 436776
rect 509775 436760 509842 436794
rect 509876 436760 510045 436794
rect 509575 436754 510045 436760
rect 509575 436720 509992 436754
rect 510026 436720 510045 436754
rect 509575 436686 509594 436720
rect 509628 436704 510045 436720
rect 509628 436686 509741 436704
rect 509575 436670 509741 436686
rect 509775 436670 509842 436704
rect 509876 436670 510045 436704
rect 509575 436664 510045 436670
rect 509575 436630 509992 436664
rect 510026 436630 510045 436664
rect 509575 436596 509594 436630
rect 509628 436614 510045 436630
rect 509628 436596 509741 436614
rect 509575 436580 509741 436596
rect 509775 436580 509842 436614
rect 509876 436580 510045 436614
rect 509575 436574 510045 436580
rect 509575 436540 509992 436574
rect 510026 436540 510045 436574
rect 509575 436506 509594 436540
rect 509628 436524 510045 436540
rect 509628 436506 509741 436524
rect 509575 436490 509741 436506
rect 509775 436490 509842 436524
rect 509876 436490 510045 436524
rect 509575 436484 510045 436490
rect 509575 436450 509992 436484
rect 510026 436450 510045 436484
rect 509575 436416 509594 436450
rect 509628 436434 510045 436450
rect 509628 436416 509741 436434
rect 509575 436400 509741 436416
rect 509775 436400 509842 436434
rect 509876 436400 510045 436434
rect 509575 436394 510045 436400
rect 509575 436360 509992 436394
rect 510026 436360 510045 436394
rect 509575 436326 509594 436360
rect 509628 436344 510045 436360
rect 509628 436326 509741 436344
rect 509575 436310 509741 436326
rect 509775 436310 509842 436344
rect 509876 436310 510045 436344
rect 509575 436304 510045 436310
rect 509575 436270 509992 436304
rect 510026 436270 510045 436304
rect 509575 436236 509594 436270
rect 509628 436254 510045 436270
rect 509628 436236 509741 436254
rect 509575 436220 509741 436236
rect 509775 436220 509842 436254
rect 509876 436220 510045 436254
rect 509575 436214 510045 436220
rect 508287 436146 508306 436180
rect 508340 436164 508757 436180
rect 508340 436146 508453 436164
rect 508287 436141 508453 436146
rect 507300 436130 508453 436141
rect 508487 436130 508554 436164
rect 508588 436141 508757 436164
rect 509575 436180 509992 436214
rect 510026 436180 510045 436214
rect 510107 436836 510801 436897
rect 510107 436802 510168 436836
rect 510202 436824 510258 436836
rect 510292 436824 510348 436836
rect 510382 436824 510438 436836
rect 510214 436802 510258 436824
rect 510314 436802 510348 436824
rect 510414 436802 510438 436824
rect 510472 436824 510528 436836
rect 510472 436802 510480 436824
rect 510107 436790 510180 436802
rect 510214 436790 510280 436802
rect 510314 436790 510380 436802
rect 510414 436790 510480 436802
rect 510514 436802 510528 436824
rect 510562 436824 510618 436836
rect 510562 436802 510580 436824
rect 510514 436790 510580 436802
rect 510614 436802 510618 436824
rect 510652 436824 510708 436836
rect 510652 436802 510680 436824
rect 510742 436802 510801 436836
rect 510614 436790 510680 436802
rect 510714 436790 510801 436802
rect 510107 436746 510801 436790
rect 510107 436712 510168 436746
rect 510202 436724 510258 436746
rect 510292 436724 510348 436746
rect 510382 436724 510438 436746
rect 510214 436712 510258 436724
rect 510314 436712 510348 436724
rect 510414 436712 510438 436724
rect 510472 436724 510528 436746
rect 510472 436712 510480 436724
rect 510107 436690 510180 436712
rect 510214 436690 510280 436712
rect 510314 436690 510380 436712
rect 510414 436690 510480 436712
rect 510514 436712 510528 436724
rect 510562 436724 510618 436746
rect 510562 436712 510580 436724
rect 510514 436690 510580 436712
rect 510614 436712 510618 436724
rect 510652 436724 510708 436746
rect 510652 436712 510680 436724
rect 510742 436712 510801 436746
rect 510614 436690 510680 436712
rect 510714 436690 510801 436712
rect 510107 436656 510801 436690
rect 510107 436622 510168 436656
rect 510202 436624 510258 436656
rect 510292 436624 510348 436656
rect 510382 436624 510438 436656
rect 510214 436622 510258 436624
rect 510314 436622 510348 436624
rect 510414 436622 510438 436624
rect 510472 436624 510528 436656
rect 510472 436622 510480 436624
rect 510107 436590 510180 436622
rect 510214 436590 510280 436622
rect 510314 436590 510380 436622
rect 510414 436590 510480 436622
rect 510514 436622 510528 436624
rect 510562 436624 510618 436656
rect 510562 436622 510580 436624
rect 510514 436590 510580 436622
rect 510614 436622 510618 436624
rect 510652 436624 510708 436656
rect 510652 436622 510680 436624
rect 510742 436622 510801 436656
rect 510614 436590 510680 436622
rect 510714 436590 510801 436622
rect 510107 436566 510801 436590
rect 510107 436532 510168 436566
rect 510202 436532 510258 436566
rect 510292 436532 510348 436566
rect 510382 436532 510438 436566
rect 510472 436532 510528 436566
rect 510562 436532 510618 436566
rect 510652 436532 510708 436566
rect 510742 436532 510801 436566
rect 510107 436524 510801 436532
rect 510107 436490 510180 436524
rect 510214 436490 510280 436524
rect 510314 436490 510380 436524
rect 510414 436490 510480 436524
rect 510514 436490 510580 436524
rect 510614 436490 510680 436524
rect 510714 436490 510801 436524
rect 510107 436476 510801 436490
rect 510107 436442 510168 436476
rect 510202 436442 510258 436476
rect 510292 436442 510348 436476
rect 510382 436442 510438 436476
rect 510472 436442 510528 436476
rect 510562 436442 510618 436476
rect 510652 436442 510708 436476
rect 510742 436442 510801 436476
rect 510107 436424 510801 436442
rect 510107 436390 510180 436424
rect 510214 436390 510280 436424
rect 510314 436390 510380 436424
rect 510414 436390 510480 436424
rect 510514 436390 510580 436424
rect 510614 436390 510680 436424
rect 510714 436390 510801 436424
rect 510107 436386 510801 436390
rect 510107 436352 510168 436386
rect 510202 436352 510258 436386
rect 510292 436352 510348 436386
rect 510382 436352 510438 436386
rect 510472 436352 510528 436386
rect 510562 436352 510618 436386
rect 510652 436352 510708 436386
rect 510742 436352 510801 436386
rect 510107 436324 510801 436352
rect 510107 436296 510180 436324
rect 510214 436296 510280 436324
rect 510314 436296 510380 436324
rect 510414 436296 510480 436324
rect 510107 436262 510168 436296
rect 510214 436290 510258 436296
rect 510314 436290 510348 436296
rect 510414 436290 510438 436296
rect 510202 436262 510258 436290
rect 510292 436262 510348 436290
rect 510382 436262 510438 436290
rect 510472 436290 510480 436296
rect 510514 436296 510580 436324
rect 510514 436290 510528 436296
rect 510472 436262 510528 436290
rect 510562 436290 510580 436296
rect 510614 436296 510680 436324
rect 510714 436296 510801 436324
rect 510614 436290 510618 436296
rect 510562 436262 510618 436290
rect 510652 436290 510680 436296
rect 510652 436262 510708 436290
rect 510742 436262 510801 436296
rect 510107 436203 510801 436262
rect 510863 436866 510882 436900
rect 510916 436884 511333 436900
rect 512151 436940 512317 436959
rect 512351 436940 512418 436974
rect 512452 436959 513605 436974
rect 512452 436940 512621 436959
rect 512151 436934 512621 436940
rect 512151 436900 512568 436934
rect 512602 436900 512621 436934
rect 510916 436866 511029 436884
rect 510863 436850 511029 436866
rect 511063 436850 511130 436884
rect 511164 436850 511333 436884
rect 510863 436844 511333 436850
rect 510863 436810 511280 436844
rect 511314 436810 511333 436844
rect 510863 436776 510882 436810
rect 510916 436794 511333 436810
rect 510916 436776 511029 436794
rect 510863 436760 511029 436776
rect 511063 436760 511130 436794
rect 511164 436760 511333 436794
rect 510863 436754 511333 436760
rect 510863 436720 511280 436754
rect 511314 436720 511333 436754
rect 510863 436686 510882 436720
rect 510916 436704 511333 436720
rect 510916 436686 511029 436704
rect 510863 436670 511029 436686
rect 511063 436670 511130 436704
rect 511164 436670 511333 436704
rect 510863 436664 511333 436670
rect 510863 436630 511280 436664
rect 511314 436630 511333 436664
rect 510863 436596 510882 436630
rect 510916 436614 511333 436630
rect 510916 436596 511029 436614
rect 510863 436580 511029 436596
rect 511063 436580 511130 436614
rect 511164 436580 511333 436614
rect 510863 436574 511333 436580
rect 510863 436540 511280 436574
rect 511314 436540 511333 436574
rect 510863 436506 510882 436540
rect 510916 436524 511333 436540
rect 510916 436506 511029 436524
rect 510863 436490 511029 436506
rect 511063 436490 511130 436524
rect 511164 436490 511333 436524
rect 510863 436484 511333 436490
rect 510863 436450 511280 436484
rect 511314 436450 511333 436484
rect 510863 436416 510882 436450
rect 510916 436434 511333 436450
rect 510916 436416 511029 436434
rect 510863 436400 511029 436416
rect 511063 436400 511130 436434
rect 511164 436400 511333 436434
rect 510863 436394 511333 436400
rect 510863 436360 511280 436394
rect 511314 436360 511333 436394
rect 510863 436326 510882 436360
rect 510916 436344 511333 436360
rect 510916 436326 511029 436344
rect 510863 436310 511029 436326
rect 511063 436310 511130 436344
rect 511164 436310 511333 436344
rect 510863 436304 511333 436310
rect 510863 436270 511280 436304
rect 511314 436270 511333 436304
rect 510863 436236 510882 436270
rect 510916 436254 511333 436270
rect 510916 436236 511029 436254
rect 510863 436220 511029 436236
rect 511063 436220 511130 436254
rect 511164 436220 511333 436254
rect 510863 436214 511333 436220
rect 509575 436146 509594 436180
rect 509628 436164 510045 436180
rect 509628 436146 509741 436164
rect 509575 436141 509741 436146
rect 508588 436130 509741 436141
rect 509775 436130 509842 436164
rect 509876 436141 510045 436164
rect 510863 436180 511280 436214
rect 511314 436180 511333 436214
rect 511395 436836 512089 436897
rect 511395 436802 511456 436836
rect 511490 436824 511546 436836
rect 511580 436824 511636 436836
rect 511670 436824 511726 436836
rect 511502 436802 511546 436824
rect 511602 436802 511636 436824
rect 511702 436802 511726 436824
rect 511760 436824 511816 436836
rect 511760 436802 511768 436824
rect 511395 436790 511468 436802
rect 511502 436790 511568 436802
rect 511602 436790 511668 436802
rect 511702 436790 511768 436802
rect 511802 436802 511816 436824
rect 511850 436824 511906 436836
rect 511850 436802 511868 436824
rect 511802 436790 511868 436802
rect 511902 436802 511906 436824
rect 511940 436824 511996 436836
rect 511940 436802 511968 436824
rect 512030 436802 512089 436836
rect 511902 436790 511968 436802
rect 512002 436790 512089 436802
rect 511395 436746 512089 436790
rect 511395 436712 511456 436746
rect 511490 436724 511546 436746
rect 511580 436724 511636 436746
rect 511670 436724 511726 436746
rect 511502 436712 511546 436724
rect 511602 436712 511636 436724
rect 511702 436712 511726 436724
rect 511760 436724 511816 436746
rect 511760 436712 511768 436724
rect 511395 436690 511468 436712
rect 511502 436690 511568 436712
rect 511602 436690 511668 436712
rect 511702 436690 511768 436712
rect 511802 436712 511816 436724
rect 511850 436724 511906 436746
rect 511850 436712 511868 436724
rect 511802 436690 511868 436712
rect 511902 436712 511906 436724
rect 511940 436724 511996 436746
rect 511940 436712 511968 436724
rect 512030 436712 512089 436746
rect 511902 436690 511968 436712
rect 512002 436690 512089 436712
rect 511395 436656 512089 436690
rect 511395 436622 511456 436656
rect 511490 436624 511546 436656
rect 511580 436624 511636 436656
rect 511670 436624 511726 436656
rect 511502 436622 511546 436624
rect 511602 436622 511636 436624
rect 511702 436622 511726 436624
rect 511760 436624 511816 436656
rect 511760 436622 511768 436624
rect 511395 436590 511468 436622
rect 511502 436590 511568 436622
rect 511602 436590 511668 436622
rect 511702 436590 511768 436622
rect 511802 436622 511816 436624
rect 511850 436624 511906 436656
rect 511850 436622 511868 436624
rect 511802 436590 511868 436622
rect 511902 436622 511906 436624
rect 511940 436624 511996 436656
rect 511940 436622 511968 436624
rect 512030 436622 512089 436656
rect 511902 436590 511968 436622
rect 512002 436590 512089 436622
rect 511395 436566 512089 436590
rect 511395 436532 511456 436566
rect 511490 436532 511546 436566
rect 511580 436532 511636 436566
rect 511670 436532 511726 436566
rect 511760 436532 511816 436566
rect 511850 436532 511906 436566
rect 511940 436532 511996 436566
rect 512030 436532 512089 436566
rect 511395 436524 512089 436532
rect 511395 436490 511468 436524
rect 511502 436490 511568 436524
rect 511602 436490 511668 436524
rect 511702 436490 511768 436524
rect 511802 436490 511868 436524
rect 511902 436490 511968 436524
rect 512002 436490 512089 436524
rect 511395 436476 512089 436490
rect 511395 436442 511456 436476
rect 511490 436442 511546 436476
rect 511580 436442 511636 436476
rect 511670 436442 511726 436476
rect 511760 436442 511816 436476
rect 511850 436442 511906 436476
rect 511940 436442 511996 436476
rect 512030 436442 512089 436476
rect 511395 436424 512089 436442
rect 511395 436390 511468 436424
rect 511502 436390 511568 436424
rect 511602 436390 511668 436424
rect 511702 436390 511768 436424
rect 511802 436390 511868 436424
rect 511902 436390 511968 436424
rect 512002 436390 512089 436424
rect 511395 436386 512089 436390
rect 511395 436352 511456 436386
rect 511490 436352 511546 436386
rect 511580 436352 511636 436386
rect 511670 436352 511726 436386
rect 511760 436352 511816 436386
rect 511850 436352 511906 436386
rect 511940 436352 511996 436386
rect 512030 436352 512089 436386
rect 511395 436324 512089 436352
rect 511395 436296 511468 436324
rect 511502 436296 511568 436324
rect 511602 436296 511668 436324
rect 511702 436296 511768 436324
rect 511395 436262 511456 436296
rect 511502 436290 511546 436296
rect 511602 436290 511636 436296
rect 511702 436290 511726 436296
rect 511490 436262 511546 436290
rect 511580 436262 511636 436290
rect 511670 436262 511726 436290
rect 511760 436290 511768 436296
rect 511802 436296 511868 436324
rect 511802 436290 511816 436296
rect 511760 436262 511816 436290
rect 511850 436290 511868 436296
rect 511902 436296 511968 436324
rect 512002 436296 512089 436324
rect 511902 436290 511906 436296
rect 511850 436262 511906 436290
rect 511940 436290 511968 436296
rect 511940 436262 511996 436290
rect 512030 436262 512089 436296
rect 511395 436203 512089 436262
rect 512151 436866 512170 436900
rect 512204 436884 512621 436900
rect 513439 436940 513605 436959
rect 513639 436940 513674 436974
rect 513439 436900 513674 436940
rect 512204 436866 512317 436884
rect 512151 436850 512317 436866
rect 512351 436850 512418 436884
rect 512452 436850 512621 436884
rect 512151 436844 512621 436850
rect 512151 436810 512568 436844
rect 512602 436810 512621 436844
rect 512151 436776 512170 436810
rect 512204 436794 512621 436810
rect 512204 436776 512317 436794
rect 512151 436760 512317 436776
rect 512351 436760 512418 436794
rect 512452 436760 512621 436794
rect 512151 436754 512621 436760
rect 512151 436720 512568 436754
rect 512602 436720 512621 436754
rect 512151 436686 512170 436720
rect 512204 436704 512621 436720
rect 512204 436686 512317 436704
rect 512151 436670 512317 436686
rect 512351 436670 512418 436704
rect 512452 436670 512621 436704
rect 512151 436664 512621 436670
rect 512151 436630 512568 436664
rect 512602 436630 512621 436664
rect 512151 436596 512170 436630
rect 512204 436614 512621 436630
rect 512204 436596 512317 436614
rect 512151 436580 512317 436596
rect 512351 436580 512418 436614
rect 512452 436580 512621 436614
rect 512151 436574 512621 436580
rect 512151 436540 512568 436574
rect 512602 436540 512621 436574
rect 512151 436506 512170 436540
rect 512204 436524 512621 436540
rect 512204 436506 512317 436524
rect 512151 436490 512317 436506
rect 512351 436490 512418 436524
rect 512452 436490 512621 436524
rect 512151 436484 512621 436490
rect 512151 436450 512568 436484
rect 512602 436450 512621 436484
rect 512151 436416 512170 436450
rect 512204 436434 512621 436450
rect 512204 436416 512317 436434
rect 512151 436400 512317 436416
rect 512351 436400 512418 436434
rect 512452 436400 512621 436434
rect 512151 436394 512621 436400
rect 512151 436360 512568 436394
rect 512602 436360 512621 436394
rect 512151 436326 512170 436360
rect 512204 436344 512621 436360
rect 512204 436326 512317 436344
rect 512151 436310 512317 436326
rect 512351 436310 512418 436344
rect 512452 436310 512621 436344
rect 512151 436304 512621 436310
rect 512151 436270 512568 436304
rect 512602 436270 512621 436304
rect 512151 436236 512170 436270
rect 512204 436254 512621 436270
rect 512204 436236 512317 436254
rect 512151 436220 512317 436236
rect 512351 436220 512418 436254
rect 512452 436220 512621 436254
rect 512151 436214 512621 436220
rect 510863 436146 510882 436180
rect 510916 436164 511333 436180
rect 510916 436146 511029 436164
rect 510863 436141 511029 436146
rect 509876 436130 511029 436141
rect 511063 436130 511130 436164
rect 511164 436141 511333 436164
rect 512151 436180 512568 436214
rect 512602 436180 512621 436214
rect 512683 436836 513377 436897
rect 512683 436802 512744 436836
rect 512778 436824 512834 436836
rect 512868 436824 512924 436836
rect 512958 436824 513014 436836
rect 512790 436802 512834 436824
rect 512890 436802 512924 436824
rect 512990 436802 513014 436824
rect 513048 436824 513104 436836
rect 513048 436802 513056 436824
rect 512683 436790 512756 436802
rect 512790 436790 512856 436802
rect 512890 436790 512956 436802
rect 512990 436790 513056 436802
rect 513090 436802 513104 436824
rect 513138 436824 513194 436836
rect 513138 436802 513156 436824
rect 513090 436790 513156 436802
rect 513190 436802 513194 436824
rect 513228 436824 513284 436836
rect 513228 436802 513256 436824
rect 513318 436802 513377 436836
rect 513190 436790 513256 436802
rect 513290 436790 513377 436802
rect 512683 436746 513377 436790
rect 512683 436712 512744 436746
rect 512778 436724 512834 436746
rect 512868 436724 512924 436746
rect 512958 436724 513014 436746
rect 512790 436712 512834 436724
rect 512890 436712 512924 436724
rect 512990 436712 513014 436724
rect 513048 436724 513104 436746
rect 513048 436712 513056 436724
rect 512683 436690 512756 436712
rect 512790 436690 512856 436712
rect 512890 436690 512956 436712
rect 512990 436690 513056 436712
rect 513090 436712 513104 436724
rect 513138 436724 513194 436746
rect 513138 436712 513156 436724
rect 513090 436690 513156 436712
rect 513190 436712 513194 436724
rect 513228 436724 513284 436746
rect 513228 436712 513256 436724
rect 513318 436712 513377 436746
rect 513190 436690 513256 436712
rect 513290 436690 513377 436712
rect 512683 436656 513377 436690
rect 512683 436622 512744 436656
rect 512778 436624 512834 436656
rect 512868 436624 512924 436656
rect 512958 436624 513014 436656
rect 512790 436622 512834 436624
rect 512890 436622 512924 436624
rect 512990 436622 513014 436624
rect 513048 436624 513104 436656
rect 513048 436622 513056 436624
rect 512683 436590 512756 436622
rect 512790 436590 512856 436622
rect 512890 436590 512956 436622
rect 512990 436590 513056 436622
rect 513090 436622 513104 436624
rect 513138 436624 513194 436656
rect 513138 436622 513156 436624
rect 513090 436590 513156 436622
rect 513190 436622 513194 436624
rect 513228 436624 513284 436656
rect 513228 436622 513256 436624
rect 513318 436622 513377 436656
rect 513190 436590 513256 436622
rect 513290 436590 513377 436622
rect 512683 436566 513377 436590
rect 512683 436532 512744 436566
rect 512778 436532 512834 436566
rect 512868 436532 512924 436566
rect 512958 436532 513014 436566
rect 513048 436532 513104 436566
rect 513138 436532 513194 436566
rect 513228 436532 513284 436566
rect 513318 436532 513377 436566
rect 512683 436524 513377 436532
rect 512683 436490 512756 436524
rect 512790 436490 512856 436524
rect 512890 436490 512956 436524
rect 512990 436490 513056 436524
rect 513090 436490 513156 436524
rect 513190 436490 513256 436524
rect 513290 436490 513377 436524
rect 512683 436476 513377 436490
rect 512683 436442 512744 436476
rect 512778 436442 512834 436476
rect 512868 436442 512924 436476
rect 512958 436442 513014 436476
rect 513048 436442 513104 436476
rect 513138 436442 513194 436476
rect 513228 436442 513284 436476
rect 513318 436442 513377 436476
rect 512683 436424 513377 436442
rect 512683 436390 512756 436424
rect 512790 436390 512856 436424
rect 512890 436390 512956 436424
rect 512990 436390 513056 436424
rect 513090 436390 513156 436424
rect 513190 436390 513256 436424
rect 513290 436390 513377 436424
rect 512683 436386 513377 436390
rect 512683 436352 512744 436386
rect 512778 436352 512834 436386
rect 512868 436352 512924 436386
rect 512958 436352 513014 436386
rect 513048 436352 513104 436386
rect 513138 436352 513194 436386
rect 513228 436352 513284 436386
rect 513318 436352 513377 436386
rect 512683 436324 513377 436352
rect 512683 436296 512756 436324
rect 512790 436296 512856 436324
rect 512890 436296 512956 436324
rect 512990 436296 513056 436324
rect 512683 436262 512744 436296
rect 512790 436290 512834 436296
rect 512890 436290 512924 436296
rect 512990 436290 513014 436296
rect 512778 436262 512834 436290
rect 512868 436262 512924 436290
rect 512958 436262 513014 436290
rect 513048 436290 513056 436296
rect 513090 436296 513156 436324
rect 513090 436290 513104 436296
rect 513048 436262 513104 436290
rect 513138 436290 513156 436296
rect 513190 436296 513256 436324
rect 513290 436296 513377 436324
rect 513190 436290 513194 436296
rect 513138 436262 513194 436290
rect 513228 436290 513256 436296
rect 513228 436262 513284 436290
rect 513318 436262 513377 436296
rect 512683 436203 513377 436262
rect 513439 436866 513458 436900
rect 513492 436884 513674 436900
rect 513492 436866 513605 436884
rect 513439 436850 513605 436866
rect 513639 436850 513674 436884
rect 513439 436810 513674 436850
rect 513439 436776 513458 436810
rect 513492 436794 513674 436810
rect 513492 436776 513605 436794
rect 513439 436760 513605 436776
rect 513639 436760 513674 436794
rect 513439 436720 513674 436760
rect 513439 436686 513458 436720
rect 513492 436704 513674 436720
rect 513492 436686 513605 436704
rect 513439 436670 513605 436686
rect 513639 436670 513674 436704
rect 513439 436630 513674 436670
rect 513439 436596 513458 436630
rect 513492 436614 513674 436630
rect 513492 436596 513605 436614
rect 513439 436580 513605 436596
rect 513639 436580 513674 436614
rect 513439 436540 513674 436580
rect 513439 436506 513458 436540
rect 513492 436524 513674 436540
rect 513492 436506 513605 436524
rect 513439 436490 513605 436506
rect 513639 436490 513674 436524
rect 513439 436450 513674 436490
rect 513439 436416 513458 436450
rect 513492 436434 513674 436450
rect 513492 436416 513605 436434
rect 513439 436400 513605 436416
rect 513639 436400 513674 436434
rect 513439 436360 513674 436400
rect 513439 436326 513458 436360
rect 513492 436344 513674 436360
rect 513492 436326 513605 436344
rect 513439 436310 513605 436326
rect 513639 436310 513674 436344
rect 513439 436270 513674 436310
rect 513439 436236 513458 436270
rect 513492 436254 513674 436270
rect 513492 436236 513605 436254
rect 513439 436220 513605 436236
rect 513639 436220 513674 436254
rect 512151 436146 512170 436180
rect 512204 436164 512621 436180
rect 512204 436146 512317 436164
rect 512151 436141 512317 436146
rect 511164 436130 512317 436141
rect 512351 436130 512418 436164
rect 512452 436141 512621 436164
rect 513439 436180 513674 436220
rect 513439 436146 513458 436180
rect 513492 436164 513674 436180
rect 513492 436146 513605 436164
rect 513439 436141 513605 436146
rect 512452 436130 513605 436141
rect 513639 436130 513674 436164
rect 503370 436122 513674 436130
rect 501368 435972 501384 436096
rect 503370 436088 503646 436122
rect 503680 436088 503736 436122
rect 503770 436088 503826 436122
rect 503860 436088 503916 436122
rect 503950 436088 504006 436122
rect 504040 436088 504096 436122
rect 504130 436088 504186 436122
rect 504220 436088 504276 436122
rect 504310 436088 504366 436122
rect 504400 436088 504934 436122
rect 504968 436088 505024 436122
rect 505058 436088 505114 436122
rect 505148 436088 505204 436122
rect 505238 436088 505294 436122
rect 505328 436088 505384 436122
rect 505418 436088 505474 436122
rect 505508 436088 505564 436122
rect 505598 436088 505654 436122
rect 505688 436088 506222 436122
rect 506256 436088 506312 436122
rect 506346 436088 506402 436122
rect 506436 436088 506492 436122
rect 506526 436088 506582 436122
rect 506616 436088 506672 436122
rect 506706 436088 506762 436122
rect 506796 436088 506852 436122
rect 506886 436088 506942 436122
rect 506976 436088 507510 436122
rect 507544 436088 507600 436122
rect 507634 436088 507690 436122
rect 507724 436088 507780 436122
rect 507814 436088 507870 436122
rect 507904 436088 507960 436122
rect 507994 436088 508050 436122
rect 508084 436088 508140 436122
rect 508174 436088 508230 436122
rect 508264 436088 508798 436122
rect 508832 436088 508888 436122
rect 508922 436088 508978 436122
rect 509012 436088 509068 436122
rect 509102 436088 509158 436122
rect 509192 436088 509248 436122
rect 509282 436088 509338 436122
rect 509372 436088 509428 436122
rect 509462 436088 509518 436122
rect 509552 436088 510086 436122
rect 510120 436088 510176 436122
rect 510210 436088 510266 436122
rect 510300 436088 510356 436122
rect 510390 436088 510446 436122
rect 510480 436088 510536 436122
rect 510570 436088 510626 436122
rect 510660 436088 510716 436122
rect 510750 436088 510806 436122
rect 510840 436088 511374 436122
rect 511408 436088 511464 436122
rect 511498 436088 511554 436122
rect 511588 436088 511644 436122
rect 511678 436088 511734 436122
rect 511768 436088 511824 436122
rect 511858 436088 511914 436122
rect 511948 436088 512004 436122
rect 512038 436088 512094 436122
rect 512128 436088 512662 436122
rect 512696 436088 512752 436122
rect 512786 436088 512842 436122
rect 512876 436088 512932 436122
rect 512966 436088 513022 436122
rect 513056 436088 513112 436122
rect 513146 436088 513202 436122
rect 513236 436088 513292 436122
rect 513326 436088 513382 436122
rect 513416 436088 513674 436122
rect 503370 436074 513674 436088
rect 503370 436040 503402 436074
rect 503436 436040 504589 436074
rect 504623 436040 504690 436074
rect 504724 436040 505877 436074
rect 505911 436040 505978 436074
rect 506012 436040 507165 436074
rect 507199 436040 507266 436074
rect 507300 436040 508453 436074
rect 508487 436040 508554 436074
rect 508588 436040 509741 436074
rect 509775 436040 509842 436074
rect 509876 436040 511029 436074
rect 511063 436040 511130 436074
rect 511164 436040 512317 436074
rect 512351 436040 512418 436074
rect 512452 436040 513605 436074
rect 513639 436040 513674 436074
rect 503370 435973 513674 436040
rect 503370 435939 503486 435973
rect 503520 435939 503576 435973
rect 503610 435939 503666 435973
rect 503700 435939 503756 435973
rect 503790 435939 503846 435973
rect 503880 435939 503936 435973
rect 503970 435939 504026 435973
rect 504060 435939 504116 435973
rect 504150 435939 504206 435973
rect 504240 435939 504296 435973
rect 504330 435939 504386 435973
rect 504420 435939 504476 435973
rect 504510 435939 504566 435973
rect 504600 435939 504774 435973
rect 504808 435939 504864 435973
rect 504898 435939 504954 435973
rect 504988 435939 505044 435973
rect 505078 435939 505134 435973
rect 505168 435939 505224 435973
rect 505258 435939 505314 435973
rect 505348 435939 505404 435973
rect 505438 435939 505494 435973
rect 505528 435939 505584 435973
rect 505618 435939 505674 435973
rect 505708 435939 505764 435973
rect 505798 435939 505854 435973
rect 505888 435939 506062 435973
rect 506096 435939 506152 435973
rect 506186 435939 506242 435973
rect 506276 435939 506332 435973
rect 506366 435939 506422 435973
rect 506456 435939 506512 435973
rect 506546 435939 506602 435973
rect 506636 435939 506692 435973
rect 506726 435939 506782 435973
rect 506816 435939 506872 435973
rect 506906 435939 506962 435973
rect 506996 435939 507052 435973
rect 507086 435939 507142 435973
rect 507176 435939 507350 435973
rect 507384 435939 507440 435973
rect 507474 435939 507530 435973
rect 507564 435939 507620 435973
rect 507654 435939 507710 435973
rect 507744 435939 507800 435973
rect 507834 435939 507890 435973
rect 507924 435939 507980 435973
rect 508014 435939 508070 435973
rect 508104 435939 508160 435973
rect 508194 435939 508250 435973
rect 508284 435939 508340 435973
rect 508374 435939 508430 435973
rect 508464 435939 508638 435973
rect 508672 435939 508728 435973
rect 508762 435939 508818 435973
rect 508852 435939 508908 435973
rect 508942 435939 508998 435973
rect 509032 435939 509088 435973
rect 509122 435939 509178 435973
rect 509212 435939 509268 435973
rect 509302 435939 509358 435973
rect 509392 435939 509448 435973
rect 509482 435939 509538 435973
rect 509572 435939 509628 435973
rect 509662 435939 509718 435973
rect 509752 435939 509926 435973
rect 509960 435939 510016 435973
rect 510050 435939 510106 435973
rect 510140 435939 510196 435973
rect 510230 435939 510286 435973
rect 510320 435939 510376 435973
rect 510410 435939 510466 435973
rect 510500 435939 510556 435973
rect 510590 435939 510646 435973
rect 510680 435939 510736 435973
rect 510770 435939 510826 435973
rect 510860 435939 510916 435973
rect 510950 435939 511006 435973
rect 511040 435939 511214 435973
rect 511248 435939 511304 435973
rect 511338 435939 511394 435973
rect 511428 435939 511484 435973
rect 511518 435939 511574 435973
rect 511608 435939 511664 435973
rect 511698 435939 511754 435973
rect 511788 435939 511844 435973
rect 511878 435939 511934 435973
rect 511968 435939 512024 435973
rect 512058 435939 512114 435973
rect 512148 435939 512204 435973
rect 512238 435939 512294 435973
rect 512328 435939 512502 435973
rect 512536 435939 512592 435973
rect 512626 435939 512682 435973
rect 512716 435939 512772 435973
rect 512806 435939 512862 435973
rect 512896 435939 512952 435973
rect 512986 435939 513042 435973
rect 513076 435939 513132 435973
rect 513166 435939 513222 435973
rect 513256 435939 513312 435973
rect 513346 435939 513402 435973
rect 513436 435939 513492 435973
rect 513526 435939 513582 435973
rect 513616 435939 513674 435973
rect 503370 435872 513674 435939
rect 501368 435748 501384 435872
rect 503370 435838 503486 435872
rect 503520 435838 503576 435872
rect 503610 435838 503666 435872
rect 503700 435838 503756 435872
rect 503790 435838 503846 435872
rect 503880 435838 503936 435872
rect 503970 435838 504026 435872
rect 504060 435838 504116 435872
rect 504150 435838 504206 435872
rect 504240 435838 504296 435872
rect 504330 435838 504386 435872
rect 504420 435838 504476 435872
rect 504510 435838 504566 435872
rect 504600 435838 504774 435872
rect 504808 435838 504864 435872
rect 504898 435838 504954 435872
rect 504988 435838 505044 435872
rect 505078 435838 505134 435872
rect 505168 435838 505224 435872
rect 505258 435838 505314 435872
rect 505348 435838 505404 435872
rect 505438 435838 505494 435872
rect 505528 435838 505584 435872
rect 505618 435838 505674 435872
rect 505708 435838 505764 435872
rect 505798 435838 505854 435872
rect 505888 435838 506062 435872
rect 506096 435838 506152 435872
rect 506186 435838 506242 435872
rect 506276 435838 506332 435872
rect 506366 435838 506422 435872
rect 506456 435838 506512 435872
rect 506546 435838 506602 435872
rect 506636 435838 506692 435872
rect 506726 435838 506782 435872
rect 506816 435838 506872 435872
rect 506906 435838 506962 435872
rect 506996 435838 507052 435872
rect 507086 435838 507142 435872
rect 507176 435838 507350 435872
rect 507384 435838 507440 435872
rect 507474 435838 507530 435872
rect 507564 435838 507620 435872
rect 507654 435838 507710 435872
rect 507744 435838 507800 435872
rect 507834 435838 507890 435872
rect 507924 435838 507980 435872
rect 508014 435838 508070 435872
rect 508104 435838 508160 435872
rect 508194 435838 508250 435872
rect 508284 435838 508340 435872
rect 508374 435838 508430 435872
rect 508464 435838 508638 435872
rect 508672 435838 508728 435872
rect 508762 435838 508818 435872
rect 508852 435838 508908 435872
rect 508942 435838 508998 435872
rect 509032 435838 509088 435872
rect 509122 435838 509178 435872
rect 509212 435838 509268 435872
rect 509302 435838 509358 435872
rect 509392 435838 509448 435872
rect 509482 435838 509538 435872
rect 509572 435838 509628 435872
rect 509662 435838 509718 435872
rect 509752 435838 509926 435872
rect 509960 435838 510016 435872
rect 510050 435838 510106 435872
rect 510140 435838 510196 435872
rect 510230 435838 510286 435872
rect 510320 435838 510376 435872
rect 510410 435838 510466 435872
rect 510500 435838 510556 435872
rect 510590 435838 510646 435872
rect 510680 435838 510736 435872
rect 510770 435838 510826 435872
rect 510860 435838 510916 435872
rect 510950 435838 511006 435872
rect 511040 435838 511214 435872
rect 511248 435838 511304 435872
rect 511338 435838 511394 435872
rect 511428 435838 511484 435872
rect 511518 435838 511574 435872
rect 511608 435838 511664 435872
rect 511698 435838 511754 435872
rect 511788 435838 511844 435872
rect 511878 435838 511934 435872
rect 511968 435838 512024 435872
rect 512058 435838 512114 435872
rect 512148 435838 512204 435872
rect 512238 435838 512294 435872
rect 512328 435838 512502 435872
rect 512536 435838 512592 435872
rect 512626 435838 512682 435872
rect 512716 435838 512772 435872
rect 512806 435838 512862 435872
rect 512896 435838 512952 435872
rect 512986 435838 513042 435872
rect 513076 435838 513132 435872
rect 513166 435838 513222 435872
rect 513256 435838 513312 435872
rect 513346 435838 513402 435872
rect 513436 435838 513492 435872
rect 513526 435838 513582 435872
rect 513616 435838 513674 435872
rect 503370 435776 513674 435838
rect 503370 435742 503402 435776
rect 503436 435742 504589 435776
rect 504623 435742 504690 435776
rect 504724 435742 505877 435776
rect 505911 435742 505978 435776
rect 506012 435742 507165 435776
rect 507199 435742 507266 435776
rect 507300 435742 508453 435776
rect 508487 435742 508554 435776
rect 508588 435742 509741 435776
rect 509775 435742 509842 435776
rect 509876 435742 511029 435776
rect 511063 435742 511130 435776
rect 511164 435742 512317 435776
rect 512351 435742 512418 435776
rect 512452 435742 513605 435776
rect 513639 435742 513674 435776
rect 503370 435724 513674 435742
rect 503370 435690 503665 435724
rect 503699 435690 503755 435724
rect 503789 435690 503845 435724
rect 503879 435690 503935 435724
rect 503969 435690 504025 435724
rect 504059 435690 504115 435724
rect 504149 435690 504205 435724
rect 504239 435690 504295 435724
rect 504329 435690 504385 435724
rect 504419 435690 504953 435724
rect 504987 435690 505043 435724
rect 505077 435690 505133 435724
rect 505167 435690 505223 435724
rect 505257 435690 505313 435724
rect 505347 435690 505403 435724
rect 505437 435690 505493 435724
rect 505527 435690 505583 435724
rect 505617 435690 505673 435724
rect 505707 435690 506241 435724
rect 506275 435690 506331 435724
rect 506365 435690 506421 435724
rect 506455 435690 506511 435724
rect 506545 435690 506601 435724
rect 506635 435690 506691 435724
rect 506725 435690 506781 435724
rect 506815 435690 506871 435724
rect 506905 435690 506961 435724
rect 506995 435690 507529 435724
rect 507563 435690 507619 435724
rect 507653 435690 507709 435724
rect 507743 435690 507799 435724
rect 507833 435690 507889 435724
rect 507923 435690 507979 435724
rect 508013 435690 508069 435724
rect 508103 435690 508159 435724
rect 508193 435690 508249 435724
rect 508283 435690 508817 435724
rect 508851 435690 508907 435724
rect 508941 435690 508997 435724
rect 509031 435690 509087 435724
rect 509121 435690 509177 435724
rect 509211 435690 509267 435724
rect 509301 435690 509357 435724
rect 509391 435690 509447 435724
rect 509481 435690 509537 435724
rect 509571 435690 510105 435724
rect 510139 435690 510195 435724
rect 510229 435690 510285 435724
rect 510319 435690 510375 435724
rect 510409 435690 510465 435724
rect 510499 435690 510555 435724
rect 510589 435690 510645 435724
rect 510679 435690 510735 435724
rect 510769 435690 510825 435724
rect 510859 435690 511393 435724
rect 511427 435690 511483 435724
rect 511517 435690 511573 435724
rect 511607 435690 511663 435724
rect 511697 435690 511753 435724
rect 511787 435690 511843 435724
rect 511877 435690 511933 435724
rect 511967 435690 512023 435724
rect 512057 435690 512113 435724
rect 512147 435690 512681 435724
rect 512715 435690 512771 435724
rect 512805 435690 512861 435724
rect 512895 435690 512951 435724
rect 512985 435690 513041 435724
rect 513075 435690 513131 435724
rect 513165 435690 513221 435724
rect 513255 435690 513311 435724
rect 513345 435690 513401 435724
rect 513435 435690 513674 435724
rect 503370 435686 513674 435690
rect 503370 435652 503402 435686
rect 503436 435671 504589 435686
rect 503436 435652 503605 435671
rect 501368 435524 501384 435648
rect 503370 435646 503605 435652
rect 503370 435612 503552 435646
rect 503586 435612 503605 435646
rect 503370 435596 503605 435612
rect 504423 435652 504589 435671
rect 504623 435652 504690 435686
rect 504724 435671 505877 435686
rect 504724 435652 504893 435671
rect 504423 435646 504893 435652
rect 504423 435612 504840 435646
rect 504874 435612 504893 435646
rect 503370 435562 503402 435596
rect 503436 435562 503605 435596
rect 503370 435556 503605 435562
rect 503370 435522 503552 435556
rect 503586 435522 503605 435556
rect 503370 435506 503605 435522
rect 503370 435472 503402 435506
rect 503436 435472 503605 435506
rect 503370 435466 503605 435472
rect 503370 435432 503552 435466
rect 503586 435432 503605 435466
rect 501368 435300 501384 435424
rect 503370 435416 503605 435432
rect 503370 435382 503402 435416
rect 503436 435382 503605 435416
rect 503370 435376 503605 435382
rect 503370 435342 503552 435376
rect 503586 435342 503605 435376
rect 503370 435326 503605 435342
rect 503370 435292 503402 435326
rect 503436 435292 503605 435326
rect 503370 435286 503605 435292
rect 503370 435252 503552 435286
rect 503586 435252 503605 435286
rect 503370 435236 503605 435252
rect 503370 435202 503402 435236
rect 503436 435202 503605 435236
rect 501368 435076 501384 435200
rect 503370 435196 503605 435202
rect 503370 435162 503552 435196
rect 503586 435162 503605 435196
rect 503370 435146 503605 435162
rect 503370 435112 503402 435146
rect 503436 435112 503605 435146
rect 503370 435106 503605 435112
rect 503370 435072 503552 435106
rect 503586 435072 503605 435106
rect 503370 435056 503605 435072
rect 503370 435022 503402 435056
rect 503436 435022 503605 435056
rect 503370 435016 503605 435022
rect 503370 434982 503552 435016
rect 503586 434982 503605 435016
rect 501368 434852 501384 434976
rect 503370 434966 503605 434982
rect 503370 434932 503402 434966
rect 503436 434932 503605 434966
rect 503370 434926 503605 434932
rect 503370 434892 503552 434926
rect 503586 434892 503605 434926
rect 503667 435548 504361 435609
rect 503667 435514 503728 435548
rect 503762 435536 503818 435548
rect 503852 435536 503908 435548
rect 503942 435536 503998 435548
rect 503774 435514 503818 435536
rect 503874 435514 503908 435536
rect 503974 435514 503998 435536
rect 504032 435536 504088 435548
rect 504032 435514 504040 435536
rect 503667 435502 503740 435514
rect 503774 435502 503840 435514
rect 503874 435502 503940 435514
rect 503974 435502 504040 435514
rect 504074 435514 504088 435536
rect 504122 435536 504178 435548
rect 504122 435514 504140 435536
rect 504074 435502 504140 435514
rect 504174 435514 504178 435536
rect 504212 435536 504268 435548
rect 504212 435514 504240 435536
rect 504302 435514 504361 435548
rect 504174 435502 504240 435514
rect 504274 435502 504361 435514
rect 503667 435458 504361 435502
rect 503667 435424 503728 435458
rect 503762 435436 503818 435458
rect 503852 435436 503908 435458
rect 503942 435436 503998 435458
rect 503774 435424 503818 435436
rect 503874 435424 503908 435436
rect 503974 435424 503998 435436
rect 504032 435436 504088 435458
rect 504032 435424 504040 435436
rect 503667 435402 503740 435424
rect 503774 435402 503840 435424
rect 503874 435402 503940 435424
rect 503974 435402 504040 435424
rect 504074 435424 504088 435436
rect 504122 435436 504178 435458
rect 504122 435424 504140 435436
rect 504074 435402 504140 435424
rect 504174 435424 504178 435436
rect 504212 435436 504268 435458
rect 504212 435424 504240 435436
rect 504302 435424 504361 435458
rect 504174 435402 504240 435424
rect 504274 435402 504361 435424
rect 503667 435368 504361 435402
rect 503667 435334 503728 435368
rect 503762 435336 503818 435368
rect 503852 435336 503908 435368
rect 503942 435336 503998 435368
rect 503774 435334 503818 435336
rect 503874 435334 503908 435336
rect 503974 435334 503998 435336
rect 504032 435336 504088 435368
rect 504032 435334 504040 435336
rect 503667 435302 503740 435334
rect 503774 435302 503840 435334
rect 503874 435302 503940 435334
rect 503974 435302 504040 435334
rect 504074 435334 504088 435336
rect 504122 435336 504178 435368
rect 504122 435334 504140 435336
rect 504074 435302 504140 435334
rect 504174 435334 504178 435336
rect 504212 435336 504268 435368
rect 504212 435334 504240 435336
rect 504302 435334 504361 435368
rect 504174 435302 504240 435334
rect 504274 435302 504361 435334
rect 503667 435278 504361 435302
rect 503667 435244 503728 435278
rect 503762 435244 503818 435278
rect 503852 435244 503908 435278
rect 503942 435244 503998 435278
rect 504032 435244 504088 435278
rect 504122 435244 504178 435278
rect 504212 435244 504268 435278
rect 504302 435244 504361 435278
rect 503667 435236 504361 435244
rect 503667 435202 503740 435236
rect 503774 435202 503840 435236
rect 503874 435202 503940 435236
rect 503974 435202 504040 435236
rect 504074 435202 504140 435236
rect 504174 435202 504240 435236
rect 504274 435202 504361 435236
rect 503667 435188 504361 435202
rect 503667 435154 503728 435188
rect 503762 435154 503818 435188
rect 503852 435154 503908 435188
rect 503942 435154 503998 435188
rect 504032 435154 504088 435188
rect 504122 435154 504178 435188
rect 504212 435154 504268 435188
rect 504302 435154 504361 435188
rect 503667 435136 504361 435154
rect 503667 435102 503740 435136
rect 503774 435102 503840 435136
rect 503874 435102 503940 435136
rect 503974 435102 504040 435136
rect 504074 435102 504140 435136
rect 504174 435102 504240 435136
rect 504274 435102 504361 435136
rect 503667 435098 504361 435102
rect 503667 435064 503728 435098
rect 503762 435064 503818 435098
rect 503852 435064 503908 435098
rect 503942 435064 503998 435098
rect 504032 435064 504088 435098
rect 504122 435064 504178 435098
rect 504212 435064 504268 435098
rect 504302 435064 504361 435098
rect 503667 435036 504361 435064
rect 503667 435008 503740 435036
rect 503774 435008 503840 435036
rect 503874 435008 503940 435036
rect 503974 435008 504040 435036
rect 503667 434974 503728 435008
rect 503774 435002 503818 435008
rect 503874 435002 503908 435008
rect 503974 435002 503998 435008
rect 503762 434974 503818 435002
rect 503852 434974 503908 435002
rect 503942 434974 503998 435002
rect 504032 435002 504040 435008
rect 504074 435008 504140 435036
rect 504074 435002 504088 435008
rect 504032 434974 504088 435002
rect 504122 435002 504140 435008
rect 504174 435008 504240 435036
rect 504274 435008 504361 435036
rect 504174 435002 504178 435008
rect 504122 434974 504178 435002
rect 504212 435002 504240 435008
rect 504212 434974 504268 435002
rect 504302 434974 504361 435008
rect 503667 434915 504361 434974
rect 504423 435578 504442 435612
rect 504476 435596 504893 435612
rect 505711 435652 505877 435671
rect 505911 435652 505978 435686
rect 506012 435671 507165 435686
rect 506012 435652 506181 435671
rect 505711 435646 506181 435652
rect 505711 435612 506128 435646
rect 506162 435612 506181 435646
rect 504476 435578 504589 435596
rect 504423 435562 504589 435578
rect 504623 435562 504690 435596
rect 504724 435562 504893 435596
rect 504423 435556 504893 435562
rect 504423 435522 504840 435556
rect 504874 435522 504893 435556
rect 504423 435488 504442 435522
rect 504476 435506 504893 435522
rect 504476 435488 504589 435506
rect 504423 435472 504589 435488
rect 504623 435472 504690 435506
rect 504724 435472 504893 435506
rect 504423 435466 504893 435472
rect 504423 435432 504840 435466
rect 504874 435432 504893 435466
rect 504423 435398 504442 435432
rect 504476 435416 504893 435432
rect 504476 435398 504589 435416
rect 504423 435382 504589 435398
rect 504623 435382 504690 435416
rect 504724 435382 504893 435416
rect 504423 435376 504893 435382
rect 504423 435342 504840 435376
rect 504874 435342 504893 435376
rect 504423 435308 504442 435342
rect 504476 435326 504893 435342
rect 504476 435308 504589 435326
rect 504423 435292 504589 435308
rect 504623 435292 504690 435326
rect 504724 435292 504893 435326
rect 504423 435286 504893 435292
rect 504423 435252 504840 435286
rect 504874 435252 504893 435286
rect 504423 435218 504442 435252
rect 504476 435236 504893 435252
rect 504476 435218 504589 435236
rect 504423 435202 504589 435218
rect 504623 435202 504690 435236
rect 504724 435202 504893 435236
rect 504423 435196 504893 435202
rect 504423 435162 504840 435196
rect 504874 435162 504893 435196
rect 504423 435128 504442 435162
rect 504476 435146 504893 435162
rect 504476 435128 504589 435146
rect 504423 435112 504589 435128
rect 504623 435112 504690 435146
rect 504724 435112 504893 435146
rect 504423 435106 504893 435112
rect 504423 435072 504840 435106
rect 504874 435072 504893 435106
rect 504423 435038 504442 435072
rect 504476 435056 504893 435072
rect 504476 435038 504589 435056
rect 504423 435022 504589 435038
rect 504623 435022 504690 435056
rect 504724 435022 504893 435056
rect 504423 435016 504893 435022
rect 504423 434982 504840 435016
rect 504874 434982 504893 435016
rect 504423 434948 504442 434982
rect 504476 434966 504893 434982
rect 504476 434948 504589 434966
rect 504423 434932 504589 434948
rect 504623 434932 504690 434966
rect 504724 434932 504893 434966
rect 504423 434926 504893 434932
rect 503370 434876 503605 434892
rect 503370 434842 503402 434876
rect 503436 434853 503605 434876
rect 504423 434892 504840 434926
rect 504874 434892 504893 434926
rect 504955 435548 505649 435609
rect 504955 435514 505016 435548
rect 505050 435536 505106 435548
rect 505140 435536 505196 435548
rect 505230 435536 505286 435548
rect 505062 435514 505106 435536
rect 505162 435514 505196 435536
rect 505262 435514 505286 435536
rect 505320 435536 505376 435548
rect 505320 435514 505328 435536
rect 504955 435502 505028 435514
rect 505062 435502 505128 435514
rect 505162 435502 505228 435514
rect 505262 435502 505328 435514
rect 505362 435514 505376 435536
rect 505410 435536 505466 435548
rect 505410 435514 505428 435536
rect 505362 435502 505428 435514
rect 505462 435514 505466 435536
rect 505500 435536 505556 435548
rect 505500 435514 505528 435536
rect 505590 435514 505649 435548
rect 505462 435502 505528 435514
rect 505562 435502 505649 435514
rect 504955 435458 505649 435502
rect 504955 435424 505016 435458
rect 505050 435436 505106 435458
rect 505140 435436 505196 435458
rect 505230 435436 505286 435458
rect 505062 435424 505106 435436
rect 505162 435424 505196 435436
rect 505262 435424 505286 435436
rect 505320 435436 505376 435458
rect 505320 435424 505328 435436
rect 504955 435402 505028 435424
rect 505062 435402 505128 435424
rect 505162 435402 505228 435424
rect 505262 435402 505328 435424
rect 505362 435424 505376 435436
rect 505410 435436 505466 435458
rect 505410 435424 505428 435436
rect 505362 435402 505428 435424
rect 505462 435424 505466 435436
rect 505500 435436 505556 435458
rect 505500 435424 505528 435436
rect 505590 435424 505649 435458
rect 505462 435402 505528 435424
rect 505562 435402 505649 435424
rect 504955 435368 505649 435402
rect 504955 435334 505016 435368
rect 505050 435336 505106 435368
rect 505140 435336 505196 435368
rect 505230 435336 505286 435368
rect 505062 435334 505106 435336
rect 505162 435334 505196 435336
rect 505262 435334 505286 435336
rect 505320 435336 505376 435368
rect 505320 435334 505328 435336
rect 504955 435302 505028 435334
rect 505062 435302 505128 435334
rect 505162 435302 505228 435334
rect 505262 435302 505328 435334
rect 505362 435334 505376 435336
rect 505410 435336 505466 435368
rect 505410 435334 505428 435336
rect 505362 435302 505428 435334
rect 505462 435334 505466 435336
rect 505500 435336 505556 435368
rect 505500 435334 505528 435336
rect 505590 435334 505649 435368
rect 505462 435302 505528 435334
rect 505562 435302 505649 435334
rect 504955 435278 505649 435302
rect 504955 435244 505016 435278
rect 505050 435244 505106 435278
rect 505140 435244 505196 435278
rect 505230 435244 505286 435278
rect 505320 435244 505376 435278
rect 505410 435244 505466 435278
rect 505500 435244 505556 435278
rect 505590 435244 505649 435278
rect 504955 435236 505649 435244
rect 504955 435202 505028 435236
rect 505062 435202 505128 435236
rect 505162 435202 505228 435236
rect 505262 435202 505328 435236
rect 505362 435202 505428 435236
rect 505462 435202 505528 435236
rect 505562 435202 505649 435236
rect 504955 435188 505649 435202
rect 504955 435154 505016 435188
rect 505050 435154 505106 435188
rect 505140 435154 505196 435188
rect 505230 435154 505286 435188
rect 505320 435154 505376 435188
rect 505410 435154 505466 435188
rect 505500 435154 505556 435188
rect 505590 435154 505649 435188
rect 504955 435136 505649 435154
rect 504955 435102 505028 435136
rect 505062 435102 505128 435136
rect 505162 435102 505228 435136
rect 505262 435102 505328 435136
rect 505362 435102 505428 435136
rect 505462 435102 505528 435136
rect 505562 435102 505649 435136
rect 504955 435098 505649 435102
rect 504955 435064 505016 435098
rect 505050 435064 505106 435098
rect 505140 435064 505196 435098
rect 505230 435064 505286 435098
rect 505320 435064 505376 435098
rect 505410 435064 505466 435098
rect 505500 435064 505556 435098
rect 505590 435064 505649 435098
rect 504955 435036 505649 435064
rect 504955 435008 505028 435036
rect 505062 435008 505128 435036
rect 505162 435008 505228 435036
rect 505262 435008 505328 435036
rect 504955 434974 505016 435008
rect 505062 435002 505106 435008
rect 505162 435002 505196 435008
rect 505262 435002 505286 435008
rect 505050 434974 505106 435002
rect 505140 434974 505196 435002
rect 505230 434974 505286 435002
rect 505320 435002 505328 435008
rect 505362 435008 505428 435036
rect 505362 435002 505376 435008
rect 505320 434974 505376 435002
rect 505410 435002 505428 435008
rect 505462 435008 505528 435036
rect 505562 435008 505649 435036
rect 505462 435002 505466 435008
rect 505410 434974 505466 435002
rect 505500 435002 505528 435008
rect 505500 434974 505556 435002
rect 505590 434974 505649 435008
rect 504955 434915 505649 434974
rect 505711 435578 505730 435612
rect 505764 435596 506181 435612
rect 506999 435652 507165 435671
rect 507199 435652 507266 435686
rect 507300 435671 508453 435686
rect 507300 435652 507469 435671
rect 506999 435646 507469 435652
rect 506999 435612 507416 435646
rect 507450 435612 507469 435646
rect 505764 435578 505877 435596
rect 505711 435562 505877 435578
rect 505911 435562 505978 435596
rect 506012 435562 506181 435596
rect 505711 435556 506181 435562
rect 505711 435522 506128 435556
rect 506162 435522 506181 435556
rect 505711 435488 505730 435522
rect 505764 435506 506181 435522
rect 505764 435488 505877 435506
rect 505711 435472 505877 435488
rect 505911 435472 505978 435506
rect 506012 435472 506181 435506
rect 505711 435466 506181 435472
rect 505711 435432 506128 435466
rect 506162 435432 506181 435466
rect 505711 435398 505730 435432
rect 505764 435416 506181 435432
rect 505764 435398 505877 435416
rect 505711 435382 505877 435398
rect 505911 435382 505978 435416
rect 506012 435382 506181 435416
rect 505711 435376 506181 435382
rect 505711 435342 506128 435376
rect 506162 435342 506181 435376
rect 505711 435308 505730 435342
rect 505764 435326 506181 435342
rect 505764 435308 505877 435326
rect 505711 435292 505877 435308
rect 505911 435292 505978 435326
rect 506012 435292 506181 435326
rect 505711 435286 506181 435292
rect 505711 435252 506128 435286
rect 506162 435252 506181 435286
rect 505711 435218 505730 435252
rect 505764 435236 506181 435252
rect 505764 435218 505877 435236
rect 505711 435202 505877 435218
rect 505911 435202 505978 435236
rect 506012 435202 506181 435236
rect 505711 435196 506181 435202
rect 505711 435162 506128 435196
rect 506162 435162 506181 435196
rect 505711 435128 505730 435162
rect 505764 435146 506181 435162
rect 505764 435128 505877 435146
rect 505711 435112 505877 435128
rect 505911 435112 505978 435146
rect 506012 435112 506181 435146
rect 505711 435106 506181 435112
rect 505711 435072 506128 435106
rect 506162 435072 506181 435106
rect 505711 435038 505730 435072
rect 505764 435056 506181 435072
rect 505764 435038 505877 435056
rect 505711 435022 505877 435038
rect 505911 435022 505978 435056
rect 506012 435022 506181 435056
rect 505711 435016 506181 435022
rect 505711 434982 506128 435016
rect 506162 434982 506181 435016
rect 505711 434948 505730 434982
rect 505764 434966 506181 434982
rect 505764 434948 505877 434966
rect 505711 434932 505877 434948
rect 505911 434932 505978 434966
rect 506012 434932 506181 434966
rect 505711 434926 506181 434932
rect 504423 434858 504442 434892
rect 504476 434876 504893 434892
rect 504476 434858 504589 434876
rect 504423 434853 504589 434858
rect 503436 434842 504589 434853
rect 504623 434842 504690 434876
rect 504724 434853 504893 434876
rect 505711 434892 506128 434926
rect 506162 434892 506181 434926
rect 506243 435548 506937 435609
rect 506243 435514 506304 435548
rect 506338 435536 506394 435548
rect 506428 435536 506484 435548
rect 506518 435536 506574 435548
rect 506350 435514 506394 435536
rect 506450 435514 506484 435536
rect 506550 435514 506574 435536
rect 506608 435536 506664 435548
rect 506608 435514 506616 435536
rect 506243 435502 506316 435514
rect 506350 435502 506416 435514
rect 506450 435502 506516 435514
rect 506550 435502 506616 435514
rect 506650 435514 506664 435536
rect 506698 435536 506754 435548
rect 506698 435514 506716 435536
rect 506650 435502 506716 435514
rect 506750 435514 506754 435536
rect 506788 435536 506844 435548
rect 506788 435514 506816 435536
rect 506878 435514 506937 435548
rect 506750 435502 506816 435514
rect 506850 435502 506937 435514
rect 506243 435458 506937 435502
rect 506243 435424 506304 435458
rect 506338 435436 506394 435458
rect 506428 435436 506484 435458
rect 506518 435436 506574 435458
rect 506350 435424 506394 435436
rect 506450 435424 506484 435436
rect 506550 435424 506574 435436
rect 506608 435436 506664 435458
rect 506608 435424 506616 435436
rect 506243 435402 506316 435424
rect 506350 435402 506416 435424
rect 506450 435402 506516 435424
rect 506550 435402 506616 435424
rect 506650 435424 506664 435436
rect 506698 435436 506754 435458
rect 506698 435424 506716 435436
rect 506650 435402 506716 435424
rect 506750 435424 506754 435436
rect 506788 435436 506844 435458
rect 506788 435424 506816 435436
rect 506878 435424 506937 435458
rect 506750 435402 506816 435424
rect 506850 435402 506937 435424
rect 506243 435368 506937 435402
rect 506243 435334 506304 435368
rect 506338 435336 506394 435368
rect 506428 435336 506484 435368
rect 506518 435336 506574 435368
rect 506350 435334 506394 435336
rect 506450 435334 506484 435336
rect 506550 435334 506574 435336
rect 506608 435336 506664 435368
rect 506608 435334 506616 435336
rect 506243 435302 506316 435334
rect 506350 435302 506416 435334
rect 506450 435302 506516 435334
rect 506550 435302 506616 435334
rect 506650 435334 506664 435336
rect 506698 435336 506754 435368
rect 506698 435334 506716 435336
rect 506650 435302 506716 435334
rect 506750 435334 506754 435336
rect 506788 435336 506844 435368
rect 506788 435334 506816 435336
rect 506878 435334 506937 435368
rect 506750 435302 506816 435334
rect 506850 435302 506937 435334
rect 506243 435278 506937 435302
rect 506243 435244 506304 435278
rect 506338 435244 506394 435278
rect 506428 435244 506484 435278
rect 506518 435244 506574 435278
rect 506608 435244 506664 435278
rect 506698 435244 506754 435278
rect 506788 435244 506844 435278
rect 506878 435244 506937 435278
rect 506243 435236 506937 435244
rect 506243 435202 506316 435236
rect 506350 435202 506416 435236
rect 506450 435202 506516 435236
rect 506550 435202 506616 435236
rect 506650 435202 506716 435236
rect 506750 435202 506816 435236
rect 506850 435202 506937 435236
rect 506243 435188 506937 435202
rect 506243 435154 506304 435188
rect 506338 435154 506394 435188
rect 506428 435154 506484 435188
rect 506518 435154 506574 435188
rect 506608 435154 506664 435188
rect 506698 435154 506754 435188
rect 506788 435154 506844 435188
rect 506878 435154 506937 435188
rect 506243 435136 506937 435154
rect 506243 435102 506316 435136
rect 506350 435102 506416 435136
rect 506450 435102 506516 435136
rect 506550 435102 506616 435136
rect 506650 435102 506716 435136
rect 506750 435102 506816 435136
rect 506850 435102 506937 435136
rect 506243 435098 506937 435102
rect 506243 435064 506304 435098
rect 506338 435064 506394 435098
rect 506428 435064 506484 435098
rect 506518 435064 506574 435098
rect 506608 435064 506664 435098
rect 506698 435064 506754 435098
rect 506788 435064 506844 435098
rect 506878 435064 506937 435098
rect 506243 435036 506937 435064
rect 506243 435008 506316 435036
rect 506350 435008 506416 435036
rect 506450 435008 506516 435036
rect 506550 435008 506616 435036
rect 506243 434974 506304 435008
rect 506350 435002 506394 435008
rect 506450 435002 506484 435008
rect 506550 435002 506574 435008
rect 506338 434974 506394 435002
rect 506428 434974 506484 435002
rect 506518 434974 506574 435002
rect 506608 435002 506616 435008
rect 506650 435008 506716 435036
rect 506650 435002 506664 435008
rect 506608 434974 506664 435002
rect 506698 435002 506716 435008
rect 506750 435008 506816 435036
rect 506850 435008 506937 435036
rect 506750 435002 506754 435008
rect 506698 434974 506754 435002
rect 506788 435002 506816 435008
rect 506788 434974 506844 435002
rect 506878 434974 506937 435008
rect 506243 434915 506937 434974
rect 506999 435578 507018 435612
rect 507052 435596 507469 435612
rect 508287 435652 508453 435671
rect 508487 435652 508554 435686
rect 508588 435671 509741 435686
rect 508588 435652 508757 435671
rect 508287 435646 508757 435652
rect 508287 435612 508704 435646
rect 508738 435612 508757 435646
rect 507052 435578 507165 435596
rect 506999 435562 507165 435578
rect 507199 435562 507266 435596
rect 507300 435562 507469 435596
rect 506999 435556 507469 435562
rect 506999 435522 507416 435556
rect 507450 435522 507469 435556
rect 506999 435488 507018 435522
rect 507052 435506 507469 435522
rect 507052 435488 507165 435506
rect 506999 435472 507165 435488
rect 507199 435472 507266 435506
rect 507300 435472 507469 435506
rect 506999 435466 507469 435472
rect 506999 435432 507416 435466
rect 507450 435432 507469 435466
rect 506999 435398 507018 435432
rect 507052 435416 507469 435432
rect 507052 435398 507165 435416
rect 506999 435382 507165 435398
rect 507199 435382 507266 435416
rect 507300 435382 507469 435416
rect 506999 435376 507469 435382
rect 506999 435342 507416 435376
rect 507450 435342 507469 435376
rect 506999 435308 507018 435342
rect 507052 435326 507469 435342
rect 507052 435308 507165 435326
rect 506999 435292 507165 435308
rect 507199 435292 507266 435326
rect 507300 435292 507469 435326
rect 506999 435286 507469 435292
rect 506999 435252 507416 435286
rect 507450 435252 507469 435286
rect 506999 435218 507018 435252
rect 507052 435236 507469 435252
rect 507052 435218 507165 435236
rect 506999 435202 507165 435218
rect 507199 435202 507266 435236
rect 507300 435202 507469 435236
rect 506999 435196 507469 435202
rect 506999 435162 507416 435196
rect 507450 435162 507469 435196
rect 506999 435128 507018 435162
rect 507052 435146 507469 435162
rect 507052 435128 507165 435146
rect 506999 435112 507165 435128
rect 507199 435112 507266 435146
rect 507300 435112 507469 435146
rect 506999 435106 507469 435112
rect 506999 435072 507416 435106
rect 507450 435072 507469 435106
rect 506999 435038 507018 435072
rect 507052 435056 507469 435072
rect 507052 435038 507165 435056
rect 506999 435022 507165 435038
rect 507199 435022 507266 435056
rect 507300 435022 507469 435056
rect 506999 435016 507469 435022
rect 506999 434982 507416 435016
rect 507450 434982 507469 435016
rect 506999 434948 507018 434982
rect 507052 434966 507469 434982
rect 507052 434948 507165 434966
rect 506999 434932 507165 434948
rect 507199 434932 507266 434966
rect 507300 434932 507469 434966
rect 506999 434926 507469 434932
rect 505711 434858 505730 434892
rect 505764 434876 506181 434892
rect 505764 434858 505877 434876
rect 505711 434853 505877 434858
rect 504724 434842 505877 434853
rect 505911 434842 505978 434876
rect 506012 434853 506181 434876
rect 506999 434892 507416 434926
rect 507450 434892 507469 434926
rect 507531 435548 508225 435609
rect 507531 435514 507592 435548
rect 507626 435536 507682 435548
rect 507716 435536 507772 435548
rect 507806 435536 507862 435548
rect 507638 435514 507682 435536
rect 507738 435514 507772 435536
rect 507838 435514 507862 435536
rect 507896 435536 507952 435548
rect 507896 435514 507904 435536
rect 507531 435502 507604 435514
rect 507638 435502 507704 435514
rect 507738 435502 507804 435514
rect 507838 435502 507904 435514
rect 507938 435514 507952 435536
rect 507986 435536 508042 435548
rect 507986 435514 508004 435536
rect 507938 435502 508004 435514
rect 508038 435514 508042 435536
rect 508076 435536 508132 435548
rect 508076 435514 508104 435536
rect 508166 435514 508225 435548
rect 508038 435502 508104 435514
rect 508138 435502 508225 435514
rect 507531 435458 508225 435502
rect 507531 435424 507592 435458
rect 507626 435436 507682 435458
rect 507716 435436 507772 435458
rect 507806 435436 507862 435458
rect 507638 435424 507682 435436
rect 507738 435424 507772 435436
rect 507838 435424 507862 435436
rect 507896 435436 507952 435458
rect 507896 435424 507904 435436
rect 507531 435402 507604 435424
rect 507638 435402 507704 435424
rect 507738 435402 507804 435424
rect 507838 435402 507904 435424
rect 507938 435424 507952 435436
rect 507986 435436 508042 435458
rect 507986 435424 508004 435436
rect 507938 435402 508004 435424
rect 508038 435424 508042 435436
rect 508076 435436 508132 435458
rect 508076 435424 508104 435436
rect 508166 435424 508225 435458
rect 508038 435402 508104 435424
rect 508138 435402 508225 435424
rect 507531 435368 508225 435402
rect 507531 435334 507592 435368
rect 507626 435336 507682 435368
rect 507716 435336 507772 435368
rect 507806 435336 507862 435368
rect 507638 435334 507682 435336
rect 507738 435334 507772 435336
rect 507838 435334 507862 435336
rect 507896 435336 507952 435368
rect 507896 435334 507904 435336
rect 507531 435302 507604 435334
rect 507638 435302 507704 435334
rect 507738 435302 507804 435334
rect 507838 435302 507904 435334
rect 507938 435334 507952 435336
rect 507986 435336 508042 435368
rect 507986 435334 508004 435336
rect 507938 435302 508004 435334
rect 508038 435334 508042 435336
rect 508076 435336 508132 435368
rect 508076 435334 508104 435336
rect 508166 435334 508225 435368
rect 508038 435302 508104 435334
rect 508138 435302 508225 435334
rect 507531 435278 508225 435302
rect 507531 435244 507592 435278
rect 507626 435244 507682 435278
rect 507716 435244 507772 435278
rect 507806 435244 507862 435278
rect 507896 435244 507952 435278
rect 507986 435244 508042 435278
rect 508076 435244 508132 435278
rect 508166 435244 508225 435278
rect 507531 435236 508225 435244
rect 507531 435202 507604 435236
rect 507638 435202 507704 435236
rect 507738 435202 507804 435236
rect 507838 435202 507904 435236
rect 507938 435202 508004 435236
rect 508038 435202 508104 435236
rect 508138 435202 508225 435236
rect 507531 435188 508225 435202
rect 507531 435154 507592 435188
rect 507626 435154 507682 435188
rect 507716 435154 507772 435188
rect 507806 435154 507862 435188
rect 507896 435154 507952 435188
rect 507986 435154 508042 435188
rect 508076 435154 508132 435188
rect 508166 435154 508225 435188
rect 507531 435136 508225 435154
rect 507531 435102 507604 435136
rect 507638 435102 507704 435136
rect 507738 435102 507804 435136
rect 507838 435102 507904 435136
rect 507938 435102 508004 435136
rect 508038 435102 508104 435136
rect 508138 435102 508225 435136
rect 507531 435098 508225 435102
rect 507531 435064 507592 435098
rect 507626 435064 507682 435098
rect 507716 435064 507772 435098
rect 507806 435064 507862 435098
rect 507896 435064 507952 435098
rect 507986 435064 508042 435098
rect 508076 435064 508132 435098
rect 508166 435064 508225 435098
rect 507531 435036 508225 435064
rect 507531 435008 507604 435036
rect 507638 435008 507704 435036
rect 507738 435008 507804 435036
rect 507838 435008 507904 435036
rect 507531 434974 507592 435008
rect 507638 435002 507682 435008
rect 507738 435002 507772 435008
rect 507838 435002 507862 435008
rect 507626 434974 507682 435002
rect 507716 434974 507772 435002
rect 507806 434974 507862 435002
rect 507896 435002 507904 435008
rect 507938 435008 508004 435036
rect 507938 435002 507952 435008
rect 507896 434974 507952 435002
rect 507986 435002 508004 435008
rect 508038 435008 508104 435036
rect 508138 435008 508225 435036
rect 508038 435002 508042 435008
rect 507986 434974 508042 435002
rect 508076 435002 508104 435008
rect 508076 434974 508132 435002
rect 508166 434974 508225 435008
rect 507531 434915 508225 434974
rect 508287 435578 508306 435612
rect 508340 435596 508757 435612
rect 509575 435652 509741 435671
rect 509775 435652 509842 435686
rect 509876 435671 511029 435686
rect 509876 435652 510045 435671
rect 509575 435646 510045 435652
rect 509575 435612 509992 435646
rect 510026 435612 510045 435646
rect 508340 435578 508453 435596
rect 508287 435562 508453 435578
rect 508487 435562 508554 435596
rect 508588 435562 508757 435596
rect 508287 435556 508757 435562
rect 508287 435522 508704 435556
rect 508738 435522 508757 435556
rect 508287 435488 508306 435522
rect 508340 435506 508757 435522
rect 508340 435488 508453 435506
rect 508287 435472 508453 435488
rect 508487 435472 508554 435506
rect 508588 435472 508757 435506
rect 508287 435466 508757 435472
rect 508287 435432 508704 435466
rect 508738 435432 508757 435466
rect 508287 435398 508306 435432
rect 508340 435416 508757 435432
rect 508340 435398 508453 435416
rect 508287 435382 508453 435398
rect 508487 435382 508554 435416
rect 508588 435382 508757 435416
rect 508287 435376 508757 435382
rect 508287 435342 508704 435376
rect 508738 435342 508757 435376
rect 508287 435308 508306 435342
rect 508340 435326 508757 435342
rect 508340 435308 508453 435326
rect 508287 435292 508453 435308
rect 508487 435292 508554 435326
rect 508588 435292 508757 435326
rect 508287 435286 508757 435292
rect 508287 435252 508704 435286
rect 508738 435252 508757 435286
rect 508287 435218 508306 435252
rect 508340 435236 508757 435252
rect 508340 435218 508453 435236
rect 508287 435202 508453 435218
rect 508487 435202 508554 435236
rect 508588 435202 508757 435236
rect 508287 435196 508757 435202
rect 508287 435162 508704 435196
rect 508738 435162 508757 435196
rect 508287 435128 508306 435162
rect 508340 435146 508757 435162
rect 508340 435128 508453 435146
rect 508287 435112 508453 435128
rect 508487 435112 508554 435146
rect 508588 435112 508757 435146
rect 508287 435106 508757 435112
rect 508287 435072 508704 435106
rect 508738 435072 508757 435106
rect 508287 435038 508306 435072
rect 508340 435056 508757 435072
rect 508340 435038 508453 435056
rect 508287 435022 508453 435038
rect 508487 435022 508554 435056
rect 508588 435022 508757 435056
rect 508287 435016 508757 435022
rect 508287 434982 508704 435016
rect 508738 434982 508757 435016
rect 508287 434948 508306 434982
rect 508340 434966 508757 434982
rect 508340 434948 508453 434966
rect 508287 434932 508453 434948
rect 508487 434932 508554 434966
rect 508588 434932 508757 434966
rect 508287 434926 508757 434932
rect 506999 434858 507018 434892
rect 507052 434876 507469 434892
rect 507052 434858 507165 434876
rect 506999 434853 507165 434858
rect 506012 434842 507165 434853
rect 507199 434842 507266 434876
rect 507300 434853 507469 434876
rect 508287 434892 508704 434926
rect 508738 434892 508757 434926
rect 508819 435548 509513 435609
rect 508819 435514 508880 435548
rect 508914 435536 508970 435548
rect 509004 435536 509060 435548
rect 509094 435536 509150 435548
rect 508926 435514 508970 435536
rect 509026 435514 509060 435536
rect 509126 435514 509150 435536
rect 509184 435536 509240 435548
rect 509184 435514 509192 435536
rect 508819 435502 508892 435514
rect 508926 435502 508992 435514
rect 509026 435502 509092 435514
rect 509126 435502 509192 435514
rect 509226 435514 509240 435536
rect 509274 435536 509330 435548
rect 509274 435514 509292 435536
rect 509226 435502 509292 435514
rect 509326 435514 509330 435536
rect 509364 435536 509420 435548
rect 509364 435514 509392 435536
rect 509454 435514 509513 435548
rect 509326 435502 509392 435514
rect 509426 435502 509513 435514
rect 508819 435458 509513 435502
rect 508819 435424 508880 435458
rect 508914 435436 508970 435458
rect 509004 435436 509060 435458
rect 509094 435436 509150 435458
rect 508926 435424 508970 435436
rect 509026 435424 509060 435436
rect 509126 435424 509150 435436
rect 509184 435436 509240 435458
rect 509184 435424 509192 435436
rect 508819 435402 508892 435424
rect 508926 435402 508992 435424
rect 509026 435402 509092 435424
rect 509126 435402 509192 435424
rect 509226 435424 509240 435436
rect 509274 435436 509330 435458
rect 509274 435424 509292 435436
rect 509226 435402 509292 435424
rect 509326 435424 509330 435436
rect 509364 435436 509420 435458
rect 509364 435424 509392 435436
rect 509454 435424 509513 435458
rect 509326 435402 509392 435424
rect 509426 435402 509513 435424
rect 508819 435368 509513 435402
rect 508819 435334 508880 435368
rect 508914 435336 508970 435368
rect 509004 435336 509060 435368
rect 509094 435336 509150 435368
rect 508926 435334 508970 435336
rect 509026 435334 509060 435336
rect 509126 435334 509150 435336
rect 509184 435336 509240 435368
rect 509184 435334 509192 435336
rect 508819 435302 508892 435334
rect 508926 435302 508992 435334
rect 509026 435302 509092 435334
rect 509126 435302 509192 435334
rect 509226 435334 509240 435336
rect 509274 435336 509330 435368
rect 509274 435334 509292 435336
rect 509226 435302 509292 435334
rect 509326 435334 509330 435336
rect 509364 435336 509420 435368
rect 509364 435334 509392 435336
rect 509454 435334 509513 435368
rect 509326 435302 509392 435334
rect 509426 435302 509513 435334
rect 508819 435278 509513 435302
rect 508819 435244 508880 435278
rect 508914 435244 508970 435278
rect 509004 435244 509060 435278
rect 509094 435244 509150 435278
rect 509184 435244 509240 435278
rect 509274 435244 509330 435278
rect 509364 435244 509420 435278
rect 509454 435244 509513 435278
rect 508819 435236 509513 435244
rect 508819 435202 508892 435236
rect 508926 435202 508992 435236
rect 509026 435202 509092 435236
rect 509126 435202 509192 435236
rect 509226 435202 509292 435236
rect 509326 435202 509392 435236
rect 509426 435202 509513 435236
rect 508819 435188 509513 435202
rect 508819 435154 508880 435188
rect 508914 435154 508970 435188
rect 509004 435154 509060 435188
rect 509094 435154 509150 435188
rect 509184 435154 509240 435188
rect 509274 435154 509330 435188
rect 509364 435154 509420 435188
rect 509454 435154 509513 435188
rect 508819 435136 509513 435154
rect 508819 435102 508892 435136
rect 508926 435102 508992 435136
rect 509026 435102 509092 435136
rect 509126 435102 509192 435136
rect 509226 435102 509292 435136
rect 509326 435102 509392 435136
rect 509426 435102 509513 435136
rect 508819 435098 509513 435102
rect 508819 435064 508880 435098
rect 508914 435064 508970 435098
rect 509004 435064 509060 435098
rect 509094 435064 509150 435098
rect 509184 435064 509240 435098
rect 509274 435064 509330 435098
rect 509364 435064 509420 435098
rect 509454 435064 509513 435098
rect 508819 435036 509513 435064
rect 508819 435008 508892 435036
rect 508926 435008 508992 435036
rect 509026 435008 509092 435036
rect 509126 435008 509192 435036
rect 508819 434974 508880 435008
rect 508926 435002 508970 435008
rect 509026 435002 509060 435008
rect 509126 435002 509150 435008
rect 508914 434974 508970 435002
rect 509004 434974 509060 435002
rect 509094 434974 509150 435002
rect 509184 435002 509192 435008
rect 509226 435008 509292 435036
rect 509226 435002 509240 435008
rect 509184 434974 509240 435002
rect 509274 435002 509292 435008
rect 509326 435008 509392 435036
rect 509426 435008 509513 435036
rect 509326 435002 509330 435008
rect 509274 434974 509330 435002
rect 509364 435002 509392 435008
rect 509364 434974 509420 435002
rect 509454 434974 509513 435008
rect 508819 434915 509513 434974
rect 509575 435578 509594 435612
rect 509628 435596 510045 435612
rect 510863 435652 511029 435671
rect 511063 435652 511130 435686
rect 511164 435671 512317 435686
rect 511164 435652 511333 435671
rect 510863 435646 511333 435652
rect 510863 435612 511280 435646
rect 511314 435612 511333 435646
rect 509628 435578 509741 435596
rect 509575 435562 509741 435578
rect 509775 435562 509842 435596
rect 509876 435562 510045 435596
rect 509575 435556 510045 435562
rect 509575 435522 509992 435556
rect 510026 435522 510045 435556
rect 509575 435488 509594 435522
rect 509628 435506 510045 435522
rect 509628 435488 509741 435506
rect 509575 435472 509741 435488
rect 509775 435472 509842 435506
rect 509876 435472 510045 435506
rect 509575 435466 510045 435472
rect 509575 435432 509992 435466
rect 510026 435432 510045 435466
rect 509575 435398 509594 435432
rect 509628 435416 510045 435432
rect 509628 435398 509741 435416
rect 509575 435382 509741 435398
rect 509775 435382 509842 435416
rect 509876 435382 510045 435416
rect 509575 435376 510045 435382
rect 509575 435342 509992 435376
rect 510026 435342 510045 435376
rect 509575 435308 509594 435342
rect 509628 435326 510045 435342
rect 509628 435308 509741 435326
rect 509575 435292 509741 435308
rect 509775 435292 509842 435326
rect 509876 435292 510045 435326
rect 509575 435286 510045 435292
rect 509575 435252 509992 435286
rect 510026 435252 510045 435286
rect 509575 435218 509594 435252
rect 509628 435236 510045 435252
rect 509628 435218 509741 435236
rect 509575 435202 509741 435218
rect 509775 435202 509842 435236
rect 509876 435202 510045 435236
rect 509575 435196 510045 435202
rect 509575 435162 509992 435196
rect 510026 435162 510045 435196
rect 509575 435128 509594 435162
rect 509628 435146 510045 435162
rect 509628 435128 509741 435146
rect 509575 435112 509741 435128
rect 509775 435112 509842 435146
rect 509876 435112 510045 435146
rect 509575 435106 510045 435112
rect 509575 435072 509992 435106
rect 510026 435072 510045 435106
rect 509575 435038 509594 435072
rect 509628 435056 510045 435072
rect 509628 435038 509741 435056
rect 509575 435022 509741 435038
rect 509775 435022 509842 435056
rect 509876 435022 510045 435056
rect 509575 435016 510045 435022
rect 509575 434982 509992 435016
rect 510026 434982 510045 435016
rect 509575 434948 509594 434982
rect 509628 434966 510045 434982
rect 509628 434948 509741 434966
rect 509575 434932 509741 434948
rect 509775 434932 509842 434966
rect 509876 434932 510045 434966
rect 509575 434926 510045 434932
rect 508287 434858 508306 434892
rect 508340 434876 508757 434892
rect 508340 434858 508453 434876
rect 508287 434853 508453 434858
rect 507300 434842 508453 434853
rect 508487 434842 508554 434876
rect 508588 434853 508757 434876
rect 509575 434892 509992 434926
rect 510026 434892 510045 434926
rect 510107 435548 510801 435609
rect 510107 435514 510168 435548
rect 510202 435536 510258 435548
rect 510292 435536 510348 435548
rect 510382 435536 510438 435548
rect 510214 435514 510258 435536
rect 510314 435514 510348 435536
rect 510414 435514 510438 435536
rect 510472 435536 510528 435548
rect 510472 435514 510480 435536
rect 510107 435502 510180 435514
rect 510214 435502 510280 435514
rect 510314 435502 510380 435514
rect 510414 435502 510480 435514
rect 510514 435514 510528 435536
rect 510562 435536 510618 435548
rect 510562 435514 510580 435536
rect 510514 435502 510580 435514
rect 510614 435514 510618 435536
rect 510652 435536 510708 435548
rect 510652 435514 510680 435536
rect 510742 435514 510801 435548
rect 510614 435502 510680 435514
rect 510714 435502 510801 435514
rect 510107 435458 510801 435502
rect 510107 435424 510168 435458
rect 510202 435436 510258 435458
rect 510292 435436 510348 435458
rect 510382 435436 510438 435458
rect 510214 435424 510258 435436
rect 510314 435424 510348 435436
rect 510414 435424 510438 435436
rect 510472 435436 510528 435458
rect 510472 435424 510480 435436
rect 510107 435402 510180 435424
rect 510214 435402 510280 435424
rect 510314 435402 510380 435424
rect 510414 435402 510480 435424
rect 510514 435424 510528 435436
rect 510562 435436 510618 435458
rect 510562 435424 510580 435436
rect 510514 435402 510580 435424
rect 510614 435424 510618 435436
rect 510652 435436 510708 435458
rect 510652 435424 510680 435436
rect 510742 435424 510801 435458
rect 510614 435402 510680 435424
rect 510714 435402 510801 435424
rect 510107 435368 510801 435402
rect 510107 435334 510168 435368
rect 510202 435336 510258 435368
rect 510292 435336 510348 435368
rect 510382 435336 510438 435368
rect 510214 435334 510258 435336
rect 510314 435334 510348 435336
rect 510414 435334 510438 435336
rect 510472 435336 510528 435368
rect 510472 435334 510480 435336
rect 510107 435302 510180 435334
rect 510214 435302 510280 435334
rect 510314 435302 510380 435334
rect 510414 435302 510480 435334
rect 510514 435334 510528 435336
rect 510562 435336 510618 435368
rect 510562 435334 510580 435336
rect 510514 435302 510580 435334
rect 510614 435334 510618 435336
rect 510652 435336 510708 435368
rect 510652 435334 510680 435336
rect 510742 435334 510801 435368
rect 510614 435302 510680 435334
rect 510714 435302 510801 435334
rect 510107 435278 510801 435302
rect 510107 435244 510168 435278
rect 510202 435244 510258 435278
rect 510292 435244 510348 435278
rect 510382 435244 510438 435278
rect 510472 435244 510528 435278
rect 510562 435244 510618 435278
rect 510652 435244 510708 435278
rect 510742 435244 510801 435278
rect 510107 435236 510801 435244
rect 510107 435202 510180 435236
rect 510214 435202 510280 435236
rect 510314 435202 510380 435236
rect 510414 435202 510480 435236
rect 510514 435202 510580 435236
rect 510614 435202 510680 435236
rect 510714 435202 510801 435236
rect 510107 435188 510801 435202
rect 510107 435154 510168 435188
rect 510202 435154 510258 435188
rect 510292 435154 510348 435188
rect 510382 435154 510438 435188
rect 510472 435154 510528 435188
rect 510562 435154 510618 435188
rect 510652 435154 510708 435188
rect 510742 435154 510801 435188
rect 510107 435136 510801 435154
rect 510107 435102 510180 435136
rect 510214 435102 510280 435136
rect 510314 435102 510380 435136
rect 510414 435102 510480 435136
rect 510514 435102 510580 435136
rect 510614 435102 510680 435136
rect 510714 435102 510801 435136
rect 510107 435098 510801 435102
rect 510107 435064 510168 435098
rect 510202 435064 510258 435098
rect 510292 435064 510348 435098
rect 510382 435064 510438 435098
rect 510472 435064 510528 435098
rect 510562 435064 510618 435098
rect 510652 435064 510708 435098
rect 510742 435064 510801 435098
rect 510107 435036 510801 435064
rect 510107 435008 510180 435036
rect 510214 435008 510280 435036
rect 510314 435008 510380 435036
rect 510414 435008 510480 435036
rect 510107 434974 510168 435008
rect 510214 435002 510258 435008
rect 510314 435002 510348 435008
rect 510414 435002 510438 435008
rect 510202 434974 510258 435002
rect 510292 434974 510348 435002
rect 510382 434974 510438 435002
rect 510472 435002 510480 435008
rect 510514 435008 510580 435036
rect 510514 435002 510528 435008
rect 510472 434974 510528 435002
rect 510562 435002 510580 435008
rect 510614 435008 510680 435036
rect 510714 435008 510801 435036
rect 510614 435002 510618 435008
rect 510562 434974 510618 435002
rect 510652 435002 510680 435008
rect 510652 434974 510708 435002
rect 510742 434974 510801 435008
rect 510107 434915 510801 434974
rect 510863 435578 510882 435612
rect 510916 435596 511333 435612
rect 512151 435652 512317 435671
rect 512351 435652 512418 435686
rect 512452 435671 513605 435686
rect 512452 435652 512621 435671
rect 512151 435646 512621 435652
rect 512151 435612 512568 435646
rect 512602 435612 512621 435646
rect 510916 435578 511029 435596
rect 510863 435562 511029 435578
rect 511063 435562 511130 435596
rect 511164 435562 511333 435596
rect 510863 435556 511333 435562
rect 510863 435522 511280 435556
rect 511314 435522 511333 435556
rect 510863 435488 510882 435522
rect 510916 435506 511333 435522
rect 510916 435488 511029 435506
rect 510863 435472 511029 435488
rect 511063 435472 511130 435506
rect 511164 435472 511333 435506
rect 510863 435466 511333 435472
rect 510863 435432 511280 435466
rect 511314 435432 511333 435466
rect 510863 435398 510882 435432
rect 510916 435416 511333 435432
rect 510916 435398 511029 435416
rect 510863 435382 511029 435398
rect 511063 435382 511130 435416
rect 511164 435382 511333 435416
rect 510863 435376 511333 435382
rect 510863 435342 511280 435376
rect 511314 435342 511333 435376
rect 510863 435308 510882 435342
rect 510916 435326 511333 435342
rect 510916 435308 511029 435326
rect 510863 435292 511029 435308
rect 511063 435292 511130 435326
rect 511164 435292 511333 435326
rect 510863 435286 511333 435292
rect 510863 435252 511280 435286
rect 511314 435252 511333 435286
rect 510863 435218 510882 435252
rect 510916 435236 511333 435252
rect 510916 435218 511029 435236
rect 510863 435202 511029 435218
rect 511063 435202 511130 435236
rect 511164 435202 511333 435236
rect 510863 435196 511333 435202
rect 510863 435162 511280 435196
rect 511314 435162 511333 435196
rect 510863 435128 510882 435162
rect 510916 435146 511333 435162
rect 510916 435128 511029 435146
rect 510863 435112 511029 435128
rect 511063 435112 511130 435146
rect 511164 435112 511333 435146
rect 510863 435106 511333 435112
rect 510863 435072 511280 435106
rect 511314 435072 511333 435106
rect 510863 435038 510882 435072
rect 510916 435056 511333 435072
rect 510916 435038 511029 435056
rect 510863 435022 511029 435038
rect 511063 435022 511130 435056
rect 511164 435022 511333 435056
rect 510863 435016 511333 435022
rect 510863 434982 511280 435016
rect 511314 434982 511333 435016
rect 510863 434948 510882 434982
rect 510916 434966 511333 434982
rect 510916 434948 511029 434966
rect 510863 434932 511029 434948
rect 511063 434932 511130 434966
rect 511164 434932 511333 434966
rect 510863 434926 511333 434932
rect 509575 434858 509594 434892
rect 509628 434876 510045 434892
rect 509628 434858 509741 434876
rect 509575 434853 509741 434858
rect 508588 434842 509741 434853
rect 509775 434842 509842 434876
rect 509876 434853 510045 434876
rect 510863 434892 511280 434926
rect 511314 434892 511333 434926
rect 511395 435548 512089 435609
rect 511395 435514 511456 435548
rect 511490 435536 511546 435548
rect 511580 435536 511636 435548
rect 511670 435536 511726 435548
rect 511502 435514 511546 435536
rect 511602 435514 511636 435536
rect 511702 435514 511726 435536
rect 511760 435536 511816 435548
rect 511760 435514 511768 435536
rect 511395 435502 511468 435514
rect 511502 435502 511568 435514
rect 511602 435502 511668 435514
rect 511702 435502 511768 435514
rect 511802 435514 511816 435536
rect 511850 435536 511906 435548
rect 511850 435514 511868 435536
rect 511802 435502 511868 435514
rect 511902 435514 511906 435536
rect 511940 435536 511996 435548
rect 511940 435514 511968 435536
rect 512030 435514 512089 435548
rect 511902 435502 511968 435514
rect 512002 435502 512089 435514
rect 511395 435458 512089 435502
rect 511395 435424 511456 435458
rect 511490 435436 511546 435458
rect 511580 435436 511636 435458
rect 511670 435436 511726 435458
rect 511502 435424 511546 435436
rect 511602 435424 511636 435436
rect 511702 435424 511726 435436
rect 511760 435436 511816 435458
rect 511760 435424 511768 435436
rect 511395 435402 511468 435424
rect 511502 435402 511568 435424
rect 511602 435402 511668 435424
rect 511702 435402 511768 435424
rect 511802 435424 511816 435436
rect 511850 435436 511906 435458
rect 511850 435424 511868 435436
rect 511802 435402 511868 435424
rect 511902 435424 511906 435436
rect 511940 435436 511996 435458
rect 511940 435424 511968 435436
rect 512030 435424 512089 435458
rect 511902 435402 511968 435424
rect 512002 435402 512089 435424
rect 511395 435368 512089 435402
rect 511395 435334 511456 435368
rect 511490 435336 511546 435368
rect 511580 435336 511636 435368
rect 511670 435336 511726 435368
rect 511502 435334 511546 435336
rect 511602 435334 511636 435336
rect 511702 435334 511726 435336
rect 511760 435336 511816 435368
rect 511760 435334 511768 435336
rect 511395 435302 511468 435334
rect 511502 435302 511568 435334
rect 511602 435302 511668 435334
rect 511702 435302 511768 435334
rect 511802 435334 511816 435336
rect 511850 435336 511906 435368
rect 511850 435334 511868 435336
rect 511802 435302 511868 435334
rect 511902 435334 511906 435336
rect 511940 435336 511996 435368
rect 511940 435334 511968 435336
rect 512030 435334 512089 435368
rect 511902 435302 511968 435334
rect 512002 435302 512089 435334
rect 511395 435278 512089 435302
rect 511395 435244 511456 435278
rect 511490 435244 511546 435278
rect 511580 435244 511636 435278
rect 511670 435244 511726 435278
rect 511760 435244 511816 435278
rect 511850 435244 511906 435278
rect 511940 435244 511996 435278
rect 512030 435244 512089 435278
rect 511395 435236 512089 435244
rect 511395 435202 511468 435236
rect 511502 435202 511568 435236
rect 511602 435202 511668 435236
rect 511702 435202 511768 435236
rect 511802 435202 511868 435236
rect 511902 435202 511968 435236
rect 512002 435202 512089 435236
rect 511395 435188 512089 435202
rect 511395 435154 511456 435188
rect 511490 435154 511546 435188
rect 511580 435154 511636 435188
rect 511670 435154 511726 435188
rect 511760 435154 511816 435188
rect 511850 435154 511906 435188
rect 511940 435154 511996 435188
rect 512030 435154 512089 435188
rect 511395 435136 512089 435154
rect 511395 435102 511468 435136
rect 511502 435102 511568 435136
rect 511602 435102 511668 435136
rect 511702 435102 511768 435136
rect 511802 435102 511868 435136
rect 511902 435102 511968 435136
rect 512002 435102 512089 435136
rect 511395 435098 512089 435102
rect 511395 435064 511456 435098
rect 511490 435064 511546 435098
rect 511580 435064 511636 435098
rect 511670 435064 511726 435098
rect 511760 435064 511816 435098
rect 511850 435064 511906 435098
rect 511940 435064 511996 435098
rect 512030 435064 512089 435098
rect 511395 435036 512089 435064
rect 511395 435008 511468 435036
rect 511502 435008 511568 435036
rect 511602 435008 511668 435036
rect 511702 435008 511768 435036
rect 511395 434974 511456 435008
rect 511502 435002 511546 435008
rect 511602 435002 511636 435008
rect 511702 435002 511726 435008
rect 511490 434974 511546 435002
rect 511580 434974 511636 435002
rect 511670 434974 511726 435002
rect 511760 435002 511768 435008
rect 511802 435008 511868 435036
rect 511802 435002 511816 435008
rect 511760 434974 511816 435002
rect 511850 435002 511868 435008
rect 511902 435008 511968 435036
rect 512002 435008 512089 435036
rect 511902 435002 511906 435008
rect 511850 434974 511906 435002
rect 511940 435002 511968 435008
rect 511940 434974 511996 435002
rect 512030 434974 512089 435008
rect 511395 434915 512089 434974
rect 512151 435578 512170 435612
rect 512204 435596 512621 435612
rect 513439 435652 513605 435671
rect 513639 435652 513674 435686
rect 513439 435612 513674 435652
rect 512204 435578 512317 435596
rect 512151 435562 512317 435578
rect 512351 435562 512418 435596
rect 512452 435562 512621 435596
rect 512151 435556 512621 435562
rect 512151 435522 512568 435556
rect 512602 435522 512621 435556
rect 512151 435488 512170 435522
rect 512204 435506 512621 435522
rect 512204 435488 512317 435506
rect 512151 435472 512317 435488
rect 512351 435472 512418 435506
rect 512452 435472 512621 435506
rect 512151 435466 512621 435472
rect 512151 435432 512568 435466
rect 512602 435432 512621 435466
rect 512151 435398 512170 435432
rect 512204 435416 512621 435432
rect 512204 435398 512317 435416
rect 512151 435382 512317 435398
rect 512351 435382 512418 435416
rect 512452 435382 512621 435416
rect 512151 435376 512621 435382
rect 512151 435342 512568 435376
rect 512602 435342 512621 435376
rect 512151 435308 512170 435342
rect 512204 435326 512621 435342
rect 512204 435308 512317 435326
rect 512151 435292 512317 435308
rect 512351 435292 512418 435326
rect 512452 435292 512621 435326
rect 512151 435286 512621 435292
rect 512151 435252 512568 435286
rect 512602 435252 512621 435286
rect 512151 435218 512170 435252
rect 512204 435236 512621 435252
rect 512204 435218 512317 435236
rect 512151 435202 512317 435218
rect 512351 435202 512418 435236
rect 512452 435202 512621 435236
rect 512151 435196 512621 435202
rect 512151 435162 512568 435196
rect 512602 435162 512621 435196
rect 512151 435128 512170 435162
rect 512204 435146 512621 435162
rect 512204 435128 512317 435146
rect 512151 435112 512317 435128
rect 512351 435112 512418 435146
rect 512452 435112 512621 435146
rect 512151 435106 512621 435112
rect 512151 435072 512568 435106
rect 512602 435072 512621 435106
rect 512151 435038 512170 435072
rect 512204 435056 512621 435072
rect 512204 435038 512317 435056
rect 512151 435022 512317 435038
rect 512351 435022 512418 435056
rect 512452 435022 512621 435056
rect 512151 435016 512621 435022
rect 512151 434982 512568 435016
rect 512602 434982 512621 435016
rect 512151 434948 512170 434982
rect 512204 434966 512621 434982
rect 512204 434948 512317 434966
rect 512151 434932 512317 434948
rect 512351 434932 512418 434966
rect 512452 434932 512621 434966
rect 512151 434926 512621 434932
rect 510863 434858 510882 434892
rect 510916 434876 511333 434892
rect 510916 434858 511029 434876
rect 510863 434853 511029 434858
rect 509876 434842 511029 434853
rect 511063 434842 511130 434876
rect 511164 434853 511333 434876
rect 512151 434892 512568 434926
rect 512602 434892 512621 434926
rect 512683 435548 513377 435609
rect 512683 435514 512744 435548
rect 512778 435536 512834 435548
rect 512868 435536 512924 435548
rect 512958 435536 513014 435548
rect 512790 435514 512834 435536
rect 512890 435514 512924 435536
rect 512990 435514 513014 435536
rect 513048 435536 513104 435548
rect 513048 435514 513056 435536
rect 512683 435502 512756 435514
rect 512790 435502 512856 435514
rect 512890 435502 512956 435514
rect 512990 435502 513056 435514
rect 513090 435514 513104 435536
rect 513138 435536 513194 435548
rect 513138 435514 513156 435536
rect 513090 435502 513156 435514
rect 513190 435514 513194 435536
rect 513228 435536 513284 435548
rect 513228 435514 513256 435536
rect 513318 435514 513377 435548
rect 513190 435502 513256 435514
rect 513290 435502 513377 435514
rect 512683 435458 513377 435502
rect 512683 435424 512744 435458
rect 512778 435436 512834 435458
rect 512868 435436 512924 435458
rect 512958 435436 513014 435458
rect 512790 435424 512834 435436
rect 512890 435424 512924 435436
rect 512990 435424 513014 435436
rect 513048 435436 513104 435458
rect 513048 435424 513056 435436
rect 512683 435402 512756 435424
rect 512790 435402 512856 435424
rect 512890 435402 512956 435424
rect 512990 435402 513056 435424
rect 513090 435424 513104 435436
rect 513138 435436 513194 435458
rect 513138 435424 513156 435436
rect 513090 435402 513156 435424
rect 513190 435424 513194 435436
rect 513228 435436 513284 435458
rect 513228 435424 513256 435436
rect 513318 435424 513377 435458
rect 513190 435402 513256 435424
rect 513290 435402 513377 435424
rect 512683 435368 513377 435402
rect 512683 435334 512744 435368
rect 512778 435336 512834 435368
rect 512868 435336 512924 435368
rect 512958 435336 513014 435368
rect 512790 435334 512834 435336
rect 512890 435334 512924 435336
rect 512990 435334 513014 435336
rect 513048 435336 513104 435368
rect 513048 435334 513056 435336
rect 512683 435302 512756 435334
rect 512790 435302 512856 435334
rect 512890 435302 512956 435334
rect 512990 435302 513056 435334
rect 513090 435334 513104 435336
rect 513138 435336 513194 435368
rect 513138 435334 513156 435336
rect 513090 435302 513156 435334
rect 513190 435334 513194 435336
rect 513228 435336 513284 435368
rect 513228 435334 513256 435336
rect 513318 435334 513377 435368
rect 513190 435302 513256 435334
rect 513290 435302 513377 435334
rect 512683 435278 513377 435302
rect 512683 435244 512744 435278
rect 512778 435244 512834 435278
rect 512868 435244 512924 435278
rect 512958 435244 513014 435278
rect 513048 435244 513104 435278
rect 513138 435244 513194 435278
rect 513228 435244 513284 435278
rect 513318 435244 513377 435278
rect 512683 435236 513377 435244
rect 512683 435202 512756 435236
rect 512790 435202 512856 435236
rect 512890 435202 512956 435236
rect 512990 435202 513056 435236
rect 513090 435202 513156 435236
rect 513190 435202 513256 435236
rect 513290 435202 513377 435236
rect 512683 435188 513377 435202
rect 512683 435154 512744 435188
rect 512778 435154 512834 435188
rect 512868 435154 512924 435188
rect 512958 435154 513014 435188
rect 513048 435154 513104 435188
rect 513138 435154 513194 435188
rect 513228 435154 513284 435188
rect 513318 435154 513377 435188
rect 512683 435136 513377 435154
rect 512683 435102 512756 435136
rect 512790 435102 512856 435136
rect 512890 435102 512956 435136
rect 512990 435102 513056 435136
rect 513090 435102 513156 435136
rect 513190 435102 513256 435136
rect 513290 435102 513377 435136
rect 512683 435098 513377 435102
rect 512683 435064 512744 435098
rect 512778 435064 512834 435098
rect 512868 435064 512924 435098
rect 512958 435064 513014 435098
rect 513048 435064 513104 435098
rect 513138 435064 513194 435098
rect 513228 435064 513284 435098
rect 513318 435064 513377 435098
rect 512683 435036 513377 435064
rect 512683 435008 512756 435036
rect 512790 435008 512856 435036
rect 512890 435008 512956 435036
rect 512990 435008 513056 435036
rect 512683 434974 512744 435008
rect 512790 435002 512834 435008
rect 512890 435002 512924 435008
rect 512990 435002 513014 435008
rect 512778 434974 512834 435002
rect 512868 434974 512924 435002
rect 512958 434974 513014 435002
rect 513048 435002 513056 435008
rect 513090 435008 513156 435036
rect 513090 435002 513104 435008
rect 513048 434974 513104 435002
rect 513138 435002 513156 435008
rect 513190 435008 513256 435036
rect 513290 435008 513377 435036
rect 513190 435002 513194 435008
rect 513138 434974 513194 435002
rect 513228 435002 513256 435008
rect 513228 434974 513284 435002
rect 513318 434974 513377 435008
rect 512683 434915 513377 434974
rect 513439 435578 513458 435612
rect 513492 435596 513674 435612
rect 513492 435578 513605 435596
rect 513439 435562 513605 435578
rect 513639 435562 513674 435596
rect 513439 435522 513674 435562
rect 513439 435488 513458 435522
rect 513492 435506 513674 435522
rect 513492 435488 513605 435506
rect 513439 435472 513605 435488
rect 513639 435472 513674 435506
rect 513439 435432 513674 435472
rect 513439 435398 513458 435432
rect 513492 435416 513674 435432
rect 513492 435398 513605 435416
rect 513439 435382 513605 435398
rect 513639 435382 513674 435416
rect 513439 435342 513674 435382
rect 513439 435308 513458 435342
rect 513492 435326 513674 435342
rect 513492 435308 513605 435326
rect 513439 435292 513605 435308
rect 513639 435292 513674 435326
rect 513439 435252 513674 435292
rect 513439 435218 513458 435252
rect 513492 435236 513674 435252
rect 513492 435218 513605 435236
rect 513439 435202 513605 435218
rect 513639 435202 513674 435236
rect 513439 435162 513674 435202
rect 513439 435128 513458 435162
rect 513492 435146 513674 435162
rect 513492 435128 513605 435146
rect 513439 435112 513605 435128
rect 513639 435112 513674 435146
rect 513439 435072 513674 435112
rect 513439 435038 513458 435072
rect 513492 435056 513674 435072
rect 513492 435038 513605 435056
rect 513439 435022 513605 435038
rect 513639 435022 513674 435056
rect 513439 434982 513674 435022
rect 513439 434948 513458 434982
rect 513492 434966 513674 434982
rect 513492 434948 513605 434966
rect 513439 434932 513605 434948
rect 513639 434932 513674 434966
rect 512151 434858 512170 434892
rect 512204 434876 512621 434892
rect 512204 434858 512317 434876
rect 512151 434853 512317 434858
rect 511164 434842 512317 434853
rect 512351 434842 512418 434876
rect 512452 434853 512621 434876
rect 513439 434892 513674 434932
rect 513439 434858 513458 434892
rect 513492 434876 513674 434892
rect 513492 434858 513605 434876
rect 513439 434853 513605 434858
rect 512452 434842 513605 434853
rect 513639 434842 513674 434876
rect 503370 434834 513674 434842
rect 503370 434800 503646 434834
rect 503680 434800 503736 434834
rect 503770 434800 503826 434834
rect 503860 434800 503916 434834
rect 503950 434800 504006 434834
rect 504040 434800 504096 434834
rect 504130 434800 504186 434834
rect 504220 434800 504276 434834
rect 504310 434800 504366 434834
rect 504400 434800 504934 434834
rect 504968 434800 505024 434834
rect 505058 434800 505114 434834
rect 505148 434800 505204 434834
rect 505238 434800 505294 434834
rect 505328 434800 505384 434834
rect 505418 434800 505474 434834
rect 505508 434800 505564 434834
rect 505598 434800 505654 434834
rect 505688 434800 506222 434834
rect 506256 434800 506312 434834
rect 506346 434800 506402 434834
rect 506436 434800 506492 434834
rect 506526 434800 506582 434834
rect 506616 434800 506672 434834
rect 506706 434800 506762 434834
rect 506796 434800 506852 434834
rect 506886 434800 506942 434834
rect 506976 434800 507510 434834
rect 507544 434800 507600 434834
rect 507634 434800 507690 434834
rect 507724 434800 507780 434834
rect 507814 434800 507870 434834
rect 507904 434800 507960 434834
rect 507994 434800 508050 434834
rect 508084 434800 508140 434834
rect 508174 434800 508230 434834
rect 508264 434800 508798 434834
rect 508832 434800 508888 434834
rect 508922 434800 508978 434834
rect 509012 434800 509068 434834
rect 509102 434800 509158 434834
rect 509192 434800 509248 434834
rect 509282 434800 509338 434834
rect 509372 434800 509428 434834
rect 509462 434800 509518 434834
rect 509552 434800 510086 434834
rect 510120 434800 510176 434834
rect 510210 434800 510266 434834
rect 510300 434800 510356 434834
rect 510390 434800 510446 434834
rect 510480 434800 510536 434834
rect 510570 434800 510626 434834
rect 510660 434800 510716 434834
rect 510750 434800 510806 434834
rect 510840 434800 511374 434834
rect 511408 434800 511464 434834
rect 511498 434800 511554 434834
rect 511588 434800 511644 434834
rect 511678 434800 511734 434834
rect 511768 434800 511824 434834
rect 511858 434800 511914 434834
rect 511948 434800 512004 434834
rect 512038 434800 512094 434834
rect 512128 434800 512662 434834
rect 512696 434800 512752 434834
rect 512786 434800 512842 434834
rect 512876 434800 512932 434834
rect 512966 434800 513022 434834
rect 513056 434800 513112 434834
rect 513146 434800 513202 434834
rect 513236 434800 513292 434834
rect 513326 434800 513382 434834
rect 513416 434800 513674 434834
rect 503370 434786 513674 434800
rect 503370 434752 503402 434786
rect 503436 434752 504589 434786
rect 504623 434752 504690 434786
rect 504724 434752 505877 434786
rect 505911 434752 505978 434786
rect 506012 434752 507165 434786
rect 507199 434752 507266 434786
rect 507300 434752 508453 434786
rect 508487 434752 508554 434786
rect 508588 434752 509741 434786
rect 509775 434752 509842 434786
rect 509876 434752 511029 434786
rect 511063 434752 511130 434786
rect 511164 434752 512317 434786
rect 512351 434752 512418 434786
rect 512452 434752 513605 434786
rect 513639 434752 513674 434786
rect 501368 434628 501384 434752
rect 503370 434685 513674 434752
rect 503370 434651 503486 434685
rect 503520 434651 503576 434685
rect 503610 434651 503666 434685
rect 503700 434651 503756 434685
rect 503790 434651 503846 434685
rect 503880 434651 503936 434685
rect 503970 434651 504026 434685
rect 504060 434651 504116 434685
rect 504150 434651 504206 434685
rect 504240 434651 504296 434685
rect 504330 434651 504386 434685
rect 504420 434651 504476 434685
rect 504510 434651 504566 434685
rect 504600 434651 504774 434685
rect 504808 434651 504864 434685
rect 504898 434651 504954 434685
rect 504988 434651 505044 434685
rect 505078 434651 505134 434685
rect 505168 434651 505224 434685
rect 505258 434651 505314 434685
rect 505348 434651 505404 434685
rect 505438 434651 505494 434685
rect 505528 434651 505584 434685
rect 505618 434651 505674 434685
rect 505708 434651 505764 434685
rect 505798 434651 505854 434685
rect 505888 434651 506062 434685
rect 506096 434651 506152 434685
rect 506186 434651 506242 434685
rect 506276 434651 506332 434685
rect 506366 434651 506422 434685
rect 506456 434651 506512 434685
rect 506546 434651 506602 434685
rect 506636 434651 506692 434685
rect 506726 434651 506782 434685
rect 506816 434651 506872 434685
rect 506906 434651 506962 434685
rect 506996 434651 507052 434685
rect 507086 434651 507142 434685
rect 507176 434651 507350 434685
rect 507384 434651 507440 434685
rect 507474 434651 507530 434685
rect 507564 434651 507620 434685
rect 507654 434651 507710 434685
rect 507744 434651 507800 434685
rect 507834 434651 507890 434685
rect 507924 434651 507980 434685
rect 508014 434651 508070 434685
rect 508104 434651 508160 434685
rect 508194 434651 508250 434685
rect 508284 434651 508340 434685
rect 508374 434651 508430 434685
rect 508464 434651 508638 434685
rect 508672 434651 508728 434685
rect 508762 434651 508818 434685
rect 508852 434651 508908 434685
rect 508942 434651 508998 434685
rect 509032 434651 509088 434685
rect 509122 434651 509178 434685
rect 509212 434651 509268 434685
rect 509302 434651 509358 434685
rect 509392 434651 509448 434685
rect 509482 434651 509538 434685
rect 509572 434651 509628 434685
rect 509662 434651 509718 434685
rect 509752 434651 509926 434685
rect 509960 434651 510016 434685
rect 510050 434651 510106 434685
rect 510140 434651 510196 434685
rect 510230 434651 510286 434685
rect 510320 434651 510376 434685
rect 510410 434651 510466 434685
rect 510500 434651 510556 434685
rect 510590 434651 510646 434685
rect 510680 434651 510736 434685
rect 510770 434651 510826 434685
rect 510860 434651 510916 434685
rect 510950 434651 511006 434685
rect 511040 434651 511214 434685
rect 511248 434651 511304 434685
rect 511338 434651 511394 434685
rect 511428 434651 511484 434685
rect 511518 434651 511574 434685
rect 511608 434651 511664 434685
rect 511698 434651 511754 434685
rect 511788 434651 511844 434685
rect 511878 434651 511934 434685
rect 511968 434651 512024 434685
rect 512058 434651 512114 434685
rect 512148 434651 512204 434685
rect 512238 434651 512294 434685
rect 512328 434651 512502 434685
rect 512536 434651 512592 434685
rect 512626 434651 512682 434685
rect 512716 434651 512772 434685
rect 512806 434651 512862 434685
rect 512896 434651 512952 434685
rect 512986 434651 513042 434685
rect 513076 434651 513132 434685
rect 513166 434651 513222 434685
rect 513256 434651 513312 434685
rect 513346 434651 513402 434685
rect 513436 434651 513492 434685
rect 513526 434651 513582 434685
rect 513616 434651 513674 434685
rect 503370 434584 513674 434651
rect 503370 434550 503486 434584
rect 503520 434550 503576 434584
rect 503610 434550 503666 434584
rect 503700 434550 503756 434584
rect 503790 434550 503846 434584
rect 503880 434550 503936 434584
rect 503970 434550 504026 434584
rect 504060 434550 504116 434584
rect 504150 434550 504206 434584
rect 504240 434550 504296 434584
rect 504330 434550 504386 434584
rect 504420 434550 504476 434584
rect 504510 434550 504566 434584
rect 504600 434550 504774 434584
rect 504808 434550 504864 434584
rect 504898 434550 504954 434584
rect 504988 434550 505044 434584
rect 505078 434550 505134 434584
rect 505168 434550 505224 434584
rect 505258 434550 505314 434584
rect 505348 434550 505404 434584
rect 505438 434550 505494 434584
rect 505528 434550 505584 434584
rect 505618 434550 505674 434584
rect 505708 434550 505764 434584
rect 505798 434550 505854 434584
rect 505888 434550 506062 434584
rect 506096 434550 506152 434584
rect 506186 434550 506242 434584
rect 506276 434550 506332 434584
rect 506366 434550 506422 434584
rect 506456 434550 506512 434584
rect 506546 434550 506602 434584
rect 506636 434550 506692 434584
rect 506726 434550 506782 434584
rect 506816 434550 506872 434584
rect 506906 434550 506962 434584
rect 506996 434550 507052 434584
rect 507086 434550 507142 434584
rect 507176 434550 507350 434584
rect 507384 434550 507440 434584
rect 507474 434550 507530 434584
rect 507564 434550 507620 434584
rect 507654 434550 507710 434584
rect 507744 434550 507800 434584
rect 507834 434550 507890 434584
rect 507924 434550 507980 434584
rect 508014 434550 508070 434584
rect 508104 434550 508160 434584
rect 508194 434550 508250 434584
rect 508284 434550 508340 434584
rect 508374 434550 508430 434584
rect 508464 434550 508638 434584
rect 508672 434550 508728 434584
rect 508762 434550 508818 434584
rect 508852 434550 508908 434584
rect 508942 434550 508998 434584
rect 509032 434550 509088 434584
rect 509122 434550 509178 434584
rect 509212 434550 509268 434584
rect 509302 434550 509358 434584
rect 509392 434550 509448 434584
rect 509482 434550 509538 434584
rect 509572 434550 509628 434584
rect 509662 434550 509718 434584
rect 509752 434550 509926 434584
rect 509960 434550 510016 434584
rect 510050 434550 510106 434584
rect 510140 434550 510196 434584
rect 510230 434550 510286 434584
rect 510320 434550 510376 434584
rect 510410 434550 510466 434584
rect 510500 434550 510556 434584
rect 510590 434550 510646 434584
rect 510680 434550 510736 434584
rect 510770 434550 510826 434584
rect 510860 434550 510916 434584
rect 510950 434550 511006 434584
rect 511040 434550 511214 434584
rect 511248 434550 511304 434584
rect 511338 434550 511394 434584
rect 511428 434550 511484 434584
rect 511518 434550 511574 434584
rect 511608 434550 511664 434584
rect 511698 434550 511754 434584
rect 511788 434550 511844 434584
rect 511878 434550 511934 434584
rect 511968 434550 512024 434584
rect 512058 434550 512114 434584
rect 512148 434550 512204 434584
rect 512238 434550 512294 434584
rect 512328 434550 512502 434584
rect 512536 434550 512592 434584
rect 512626 434550 512682 434584
rect 512716 434550 512772 434584
rect 512806 434550 512862 434584
rect 512896 434550 512952 434584
rect 512986 434550 513042 434584
rect 513076 434550 513132 434584
rect 513166 434550 513222 434584
rect 513256 434550 513312 434584
rect 513346 434550 513402 434584
rect 513436 434550 513492 434584
rect 513526 434550 513582 434584
rect 513616 434550 513674 434584
rect 501368 434404 501384 434528
rect 503370 434488 513674 434550
rect 503370 434454 503402 434488
rect 503436 434454 504589 434488
rect 504623 434454 504690 434488
rect 504724 434454 505877 434488
rect 505911 434454 505978 434488
rect 506012 434454 507165 434488
rect 507199 434454 507266 434488
rect 507300 434454 508453 434488
rect 508487 434454 508554 434488
rect 508588 434454 509741 434488
rect 509775 434454 509842 434488
rect 509876 434454 511029 434488
rect 511063 434454 511130 434488
rect 511164 434454 512317 434488
rect 512351 434454 512418 434488
rect 512452 434454 513605 434488
rect 513639 434454 513674 434488
rect 503370 434436 513674 434454
rect 503370 434402 503665 434436
rect 503699 434402 503755 434436
rect 503789 434402 503845 434436
rect 503879 434402 503935 434436
rect 503969 434402 504025 434436
rect 504059 434402 504115 434436
rect 504149 434402 504205 434436
rect 504239 434402 504295 434436
rect 504329 434402 504385 434436
rect 504419 434402 504953 434436
rect 504987 434402 505043 434436
rect 505077 434402 505133 434436
rect 505167 434402 505223 434436
rect 505257 434402 505313 434436
rect 505347 434402 505403 434436
rect 505437 434402 505493 434436
rect 505527 434402 505583 434436
rect 505617 434402 505673 434436
rect 505707 434402 506241 434436
rect 506275 434402 506331 434436
rect 506365 434402 506421 434436
rect 506455 434402 506511 434436
rect 506545 434402 506601 434436
rect 506635 434402 506691 434436
rect 506725 434402 506781 434436
rect 506815 434402 506871 434436
rect 506905 434402 506961 434436
rect 506995 434402 507529 434436
rect 507563 434402 507619 434436
rect 507653 434402 507709 434436
rect 507743 434402 507799 434436
rect 507833 434402 507889 434436
rect 507923 434402 507979 434436
rect 508013 434402 508069 434436
rect 508103 434402 508159 434436
rect 508193 434402 508249 434436
rect 508283 434402 508817 434436
rect 508851 434402 508907 434436
rect 508941 434402 508997 434436
rect 509031 434402 509087 434436
rect 509121 434402 509177 434436
rect 509211 434402 509267 434436
rect 509301 434402 509357 434436
rect 509391 434402 509447 434436
rect 509481 434402 509537 434436
rect 509571 434402 510105 434436
rect 510139 434402 510195 434436
rect 510229 434402 510285 434436
rect 510319 434402 510375 434436
rect 510409 434402 510465 434436
rect 510499 434402 510555 434436
rect 510589 434402 510645 434436
rect 510679 434402 510735 434436
rect 510769 434402 510825 434436
rect 510859 434402 511393 434436
rect 511427 434402 511483 434436
rect 511517 434402 511573 434436
rect 511607 434402 511663 434436
rect 511697 434402 511753 434436
rect 511787 434402 511843 434436
rect 511877 434402 511933 434436
rect 511967 434402 512023 434436
rect 512057 434402 512113 434436
rect 512147 434402 512681 434436
rect 512715 434402 512771 434436
rect 512805 434402 512861 434436
rect 512895 434402 512951 434436
rect 512985 434402 513041 434436
rect 513075 434402 513131 434436
rect 513165 434402 513221 434436
rect 513255 434402 513311 434436
rect 513345 434402 513401 434436
rect 513435 434402 513674 434436
rect 503370 434398 513674 434402
rect 503370 434364 503402 434398
rect 503436 434383 504589 434398
rect 503436 434364 503605 434383
rect 503370 434358 503605 434364
rect 503370 434324 503552 434358
rect 503586 434324 503605 434358
rect 503370 434308 503605 434324
rect 504423 434364 504589 434383
rect 504623 434364 504690 434398
rect 504724 434383 505877 434398
rect 504724 434364 504893 434383
rect 504423 434358 504893 434364
rect 504423 434324 504840 434358
rect 504874 434324 504893 434358
rect 501368 434180 501384 434304
rect 503370 434274 503402 434308
rect 503436 434274 503605 434308
rect 503370 434268 503605 434274
rect 503370 434234 503552 434268
rect 503586 434234 503605 434268
rect 503370 434218 503605 434234
rect 503370 434184 503402 434218
rect 503436 434184 503605 434218
rect 503370 434178 503605 434184
rect 503370 434144 503552 434178
rect 503586 434144 503605 434178
rect 503370 434128 503605 434144
rect 503370 434094 503402 434128
rect 503436 434094 503605 434128
rect 503370 434088 503605 434094
rect 501368 433956 501384 434080
rect 503370 434054 503552 434088
rect 503586 434054 503605 434088
rect 503370 434038 503605 434054
rect 503370 434004 503402 434038
rect 503436 434004 503605 434038
rect 503370 433998 503605 434004
rect 503370 433964 503552 433998
rect 503586 433964 503605 433998
rect 503370 433948 503605 433964
rect 503370 433914 503402 433948
rect 503436 433914 503605 433948
rect 503370 433908 503605 433914
rect 503370 433874 503552 433908
rect 503586 433874 503605 433908
rect 503370 433858 503605 433874
rect 501368 433732 501384 433856
rect 503370 433824 503402 433858
rect 503436 433824 503605 433858
rect 503370 433818 503605 433824
rect 503370 433784 503552 433818
rect 503586 433784 503605 433818
rect 503370 433768 503605 433784
rect 503370 433734 503402 433768
rect 503436 433734 503605 433768
rect 503370 433728 503605 433734
rect 503370 433694 503552 433728
rect 503586 433694 503605 433728
rect 503370 433678 503605 433694
rect 503370 433644 503402 433678
rect 503436 433644 503605 433678
rect 503370 433638 503605 433644
rect 501368 433508 501384 433632
rect 503370 433604 503552 433638
rect 503586 433604 503605 433638
rect 503667 434260 504361 434321
rect 503667 434226 503728 434260
rect 503762 434248 503818 434260
rect 503852 434248 503908 434260
rect 503942 434248 503998 434260
rect 503774 434226 503818 434248
rect 503874 434226 503908 434248
rect 503974 434226 503998 434248
rect 504032 434248 504088 434260
rect 504032 434226 504040 434248
rect 503667 434214 503740 434226
rect 503774 434214 503840 434226
rect 503874 434214 503940 434226
rect 503974 434214 504040 434226
rect 504074 434226 504088 434248
rect 504122 434248 504178 434260
rect 504122 434226 504140 434248
rect 504074 434214 504140 434226
rect 504174 434226 504178 434248
rect 504212 434248 504268 434260
rect 504212 434226 504240 434248
rect 504302 434226 504361 434260
rect 504174 434214 504240 434226
rect 504274 434214 504361 434226
rect 503667 434170 504361 434214
rect 503667 434136 503728 434170
rect 503762 434148 503818 434170
rect 503852 434148 503908 434170
rect 503942 434148 503998 434170
rect 503774 434136 503818 434148
rect 503874 434136 503908 434148
rect 503974 434136 503998 434148
rect 504032 434148 504088 434170
rect 504032 434136 504040 434148
rect 503667 434114 503740 434136
rect 503774 434114 503840 434136
rect 503874 434114 503940 434136
rect 503974 434114 504040 434136
rect 504074 434136 504088 434148
rect 504122 434148 504178 434170
rect 504122 434136 504140 434148
rect 504074 434114 504140 434136
rect 504174 434136 504178 434148
rect 504212 434148 504268 434170
rect 504212 434136 504240 434148
rect 504302 434136 504361 434170
rect 504174 434114 504240 434136
rect 504274 434114 504361 434136
rect 503667 434080 504361 434114
rect 503667 434046 503728 434080
rect 503762 434048 503818 434080
rect 503852 434048 503908 434080
rect 503942 434048 503998 434080
rect 503774 434046 503818 434048
rect 503874 434046 503908 434048
rect 503974 434046 503998 434048
rect 504032 434048 504088 434080
rect 504032 434046 504040 434048
rect 503667 434014 503740 434046
rect 503774 434014 503840 434046
rect 503874 434014 503940 434046
rect 503974 434014 504040 434046
rect 504074 434046 504088 434048
rect 504122 434048 504178 434080
rect 504122 434046 504140 434048
rect 504074 434014 504140 434046
rect 504174 434046 504178 434048
rect 504212 434048 504268 434080
rect 504212 434046 504240 434048
rect 504302 434046 504361 434080
rect 504174 434014 504240 434046
rect 504274 434014 504361 434046
rect 503667 433990 504361 434014
rect 503667 433956 503728 433990
rect 503762 433956 503818 433990
rect 503852 433956 503908 433990
rect 503942 433956 503998 433990
rect 504032 433956 504088 433990
rect 504122 433956 504178 433990
rect 504212 433956 504268 433990
rect 504302 433956 504361 433990
rect 503667 433948 504361 433956
rect 503667 433914 503740 433948
rect 503774 433914 503840 433948
rect 503874 433914 503940 433948
rect 503974 433914 504040 433948
rect 504074 433914 504140 433948
rect 504174 433914 504240 433948
rect 504274 433914 504361 433948
rect 503667 433900 504361 433914
rect 503667 433866 503728 433900
rect 503762 433866 503818 433900
rect 503852 433866 503908 433900
rect 503942 433866 503998 433900
rect 504032 433866 504088 433900
rect 504122 433866 504178 433900
rect 504212 433866 504268 433900
rect 504302 433866 504361 433900
rect 503667 433848 504361 433866
rect 503667 433814 503740 433848
rect 503774 433814 503840 433848
rect 503874 433814 503940 433848
rect 503974 433814 504040 433848
rect 504074 433814 504140 433848
rect 504174 433814 504240 433848
rect 504274 433814 504361 433848
rect 503667 433810 504361 433814
rect 503667 433776 503728 433810
rect 503762 433776 503818 433810
rect 503852 433776 503908 433810
rect 503942 433776 503998 433810
rect 504032 433776 504088 433810
rect 504122 433776 504178 433810
rect 504212 433776 504268 433810
rect 504302 433776 504361 433810
rect 503667 433748 504361 433776
rect 503667 433720 503740 433748
rect 503774 433720 503840 433748
rect 503874 433720 503940 433748
rect 503974 433720 504040 433748
rect 503667 433686 503728 433720
rect 503774 433714 503818 433720
rect 503874 433714 503908 433720
rect 503974 433714 503998 433720
rect 503762 433686 503818 433714
rect 503852 433686 503908 433714
rect 503942 433686 503998 433714
rect 504032 433714 504040 433720
rect 504074 433720 504140 433748
rect 504074 433714 504088 433720
rect 504032 433686 504088 433714
rect 504122 433714 504140 433720
rect 504174 433720 504240 433748
rect 504274 433720 504361 433748
rect 504174 433714 504178 433720
rect 504122 433686 504178 433714
rect 504212 433714 504240 433720
rect 504212 433686 504268 433714
rect 504302 433686 504361 433720
rect 503667 433627 504361 433686
rect 504423 434290 504442 434324
rect 504476 434308 504893 434324
rect 505711 434364 505877 434383
rect 505911 434364 505978 434398
rect 506012 434383 507165 434398
rect 506012 434364 506181 434383
rect 505711 434358 506181 434364
rect 505711 434324 506128 434358
rect 506162 434324 506181 434358
rect 504476 434290 504589 434308
rect 504423 434274 504589 434290
rect 504623 434274 504690 434308
rect 504724 434274 504893 434308
rect 504423 434268 504893 434274
rect 504423 434234 504840 434268
rect 504874 434234 504893 434268
rect 504423 434200 504442 434234
rect 504476 434218 504893 434234
rect 504476 434200 504589 434218
rect 504423 434184 504589 434200
rect 504623 434184 504690 434218
rect 504724 434184 504893 434218
rect 504423 434178 504893 434184
rect 504423 434144 504840 434178
rect 504874 434144 504893 434178
rect 504423 434110 504442 434144
rect 504476 434128 504893 434144
rect 504476 434110 504589 434128
rect 504423 434094 504589 434110
rect 504623 434094 504690 434128
rect 504724 434094 504893 434128
rect 504423 434088 504893 434094
rect 504423 434054 504840 434088
rect 504874 434054 504893 434088
rect 504423 434020 504442 434054
rect 504476 434038 504893 434054
rect 504476 434020 504589 434038
rect 504423 434004 504589 434020
rect 504623 434004 504690 434038
rect 504724 434004 504893 434038
rect 504423 433998 504893 434004
rect 504423 433964 504840 433998
rect 504874 433964 504893 433998
rect 504423 433930 504442 433964
rect 504476 433948 504893 433964
rect 504476 433930 504589 433948
rect 504423 433914 504589 433930
rect 504623 433914 504690 433948
rect 504724 433914 504893 433948
rect 504423 433908 504893 433914
rect 504423 433874 504840 433908
rect 504874 433874 504893 433908
rect 504423 433840 504442 433874
rect 504476 433858 504893 433874
rect 504476 433840 504589 433858
rect 504423 433824 504589 433840
rect 504623 433824 504690 433858
rect 504724 433824 504893 433858
rect 504423 433818 504893 433824
rect 504423 433784 504840 433818
rect 504874 433784 504893 433818
rect 504423 433750 504442 433784
rect 504476 433768 504893 433784
rect 504476 433750 504589 433768
rect 504423 433734 504589 433750
rect 504623 433734 504690 433768
rect 504724 433734 504893 433768
rect 504423 433728 504893 433734
rect 504423 433694 504840 433728
rect 504874 433694 504893 433728
rect 504423 433660 504442 433694
rect 504476 433678 504893 433694
rect 504476 433660 504589 433678
rect 504423 433644 504589 433660
rect 504623 433644 504690 433678
rect 504724 433644 504893 433678
rect 504423 433638 504893 433644
rect 503370 433588 503605 433604
rect 503370 433554 503402 433588
rect 503436 433565 503605 433588
rect 504423 433604 504840 433638
rect 504874 433604 504893 433638
rect 504955 434260 505649 434321
rect 504955 434226 505016 434260
rect 505050 434248 505106 434260
rect 505140 434248 505196 434260
rect 505230 434248 505286 434260
rect 505062 434226 505106 434248
rect 505162 434226 505196 434248
rect 505262 434226 505286 434248
rect 505320 434248 505376 434260
rect 505320 434226 505328 434248
rect 504955 434214 505028 434226
rect 505062 434214 505128 434226
rect 505162 434214 505228 434226
rect 505262 434214 505328 434226
rect 505362 434226 505376 434248
rect 505410 434248 505466 434260
rect 505410 434226 505428 434248
rect 505362 434214 505428 434226
rect 505462 434226 505466 434248
rect 505500 434248 505556 434260
rect 505500 434226 505528 434248
rect 505590 434226 505649 434260
rect 505462 434214 505528 434226
rect 505562 434214 505649 434226
rect 504955 434170 505649 434214
rect 504955 434136 505016 434170
rect 505050 434148 505106 434170
rect 505140 434148 505196 434170
rect 505230 434148 505286 434170
rect 505062 434136 505106 434148
rect 505162 434136 505196 434148
rect 505262 434136 505286 434148
rect 505320 434148 505376 434170
rect 505320 434136 505328 434148
rect 504955 434114 505028 434136
rect 505062 434114 505128 434136
rect 505162 434114 505228 434136
rect 505262 434114 505328 434136
rect 505362 434136 505376 434148
rect 505410 434148 505466 434170
rect 505410 434136 505428 434148
rect 505362 434114 505428 434136
rect 505462 434136 505466 434148
rect 505500 434148 505556 434170
rect 505500 434136 505528 434148
rect 505590 434136 505649 434170
rect 505462 434114 505528 434136
rect 505562 434114 505649 434136
rect 504955 434080 505649 434114
rect 504955 434046 505016 434080
rect 505050 434048 505106 434080
rect 505140 434048 505196 434080
rect 505230 434048 505286 434080
rect 505062 434046 505106 434048
rect 505162 434046 505196 434048
rect 505262 434046 505286 434048
rect 505320 434048 505376 434080
rect 505320 434046 505328 434048
rect 504955 434014 505028 434046
rect 505062 434014 505128 434046
rect 505162 434014 505228 434046
rect 505262 434014 505328 434046
rect 505362 434046 505376 434048
rect 505410 434048 505466 434080
rect 505410 434046 505428 434048
rect 505362 434014 505428 434046
rect 505462 434046 505466 434048
rect 505500 434048 505556 434080
rect 505500 434046 505528 434048
rect 505590 434046 505649 434080
rect 505462 434014 505528 434046
rect 505562 434014 505649 434046
rect 504955 433990 505649 434014
rect 504955 433956 505016 433990
rect 505050 433956 505106 433990
rect 505140 433956 505196 433990
rect 505230 433956 505286 433990
rect 505320 433956 505376 433990
rect 505410 433956 505466 433990
rect 505500 433956 505556 433990
rect 505590 433956 505649 433990
rect 504955 433948 505649 433956
rect 504955 433914 505028 433948
rect 505062 433914 505128 433948
rect 505162 433914 505228 433948
rect 505262 433914 505328 433948
rect 505362 433914 505428 433948
rect 505462 433914 505528 433948
rect 505562 433914 505649 433948
rect 504955 433900 505649 433914
rect 504955 433866 505016 433900
rect 505050 433866 505106 433900
rect 505140 433866 505196 433900
rect 505230 433866 505286 433900
rect 505320 433866 505376 433900
rect 505410 433866 505466 433900
rect 505500 433866 505556 433900
rect 505590 433866 505649 433900
rect 504955 433848 505649 433866
rect 504955 433814 505028 433848
rect 505062 433814 505128 433848
rect 505162 433814 505228 433848
rect 505262 433814 505328 433848
rect 505362 433814 505428 433848
rect 505462 433814 505528 433848
rect 505562 433814 505649 433848
rect 504955 433810 505649 433814
rect 504955 433776 505016 433810
rect 505050 433776 505106 433810
rect 505140 433776 505196 433810
rect 505230 433776 505286 433810
rect 505320 433776 505376 433810
rect 505410 433776 505466 433810
rect 505500 433776 505556 433810
rect 505590 433776 505649 433810
rect 504955 433748 505649 433776
rect 504955 433720 505028 433748
rect 505062 433720 505128 433748
rect 505162 433720 505228 433748
rect 505262 433720 505328 433748
rect 504955 433686 505016 433720
rect 505062 433714 505106 433720
rect 505162 433714 505196 433720
rect 505262 433714 505286 433720
rect 505050 433686 505106 433714
rect 505140 433686 505196 433714
rect 505230 433686 505286 433714
rect 505320 433714 505328 433720
rect 505362 433720 505428 433748
rect 505362 433714 505376 433720
rect 505320 433686 505376 433714
rect 505410 433714 505428 433720
rect 505462 433720 505528 433748
rect 505562 433720 505649 433748
rect 505462 433714 505466 433720
rect 505410 433686 505466 433714
rect 505500 433714 505528 433720
rect 505500 433686 505556 433714
rect 505590 433686 505649 433720
rect 504955 433627 505649 433686
rect 505711 434290 505730 434324
rect 505764 434308 506181 434324
rect 506999 434364 507165 434383
rect 507199 434364 507266 434398
rect 507300 434383 508453 434398
rect 507300 434364 507469 434383
rect 506999 434358 507469 434364
rect 506999 434324 507416 434358
rect 507450 434324 507469 434358
rect 505764 434290 505877 434308
rect 505711 434274 505877 434290
rect 505911 434274 505978 434308
rect 506012 434274 506181 434308
rect 505711 434268 506181 434274
rect 505711 434234 506128 434268
rect 506162 434234 506181 434268
rect 505711 434200 505730 434234
rect 505764 434218 506181 434234
rect 505764 434200 505877 434218
rect 505711 434184 505877 434200
rect 505911 434184 505978 434218
rect 506012 434184 506181 434218
rect 505711 434178 506181 434184
rect 505711 434144 506128 434178
rect 506162 434144 506181 434178
rect 505711 434110 505730 434144
rect 505764 434128 506181 434144
rect 505764 434110 505877 434128
rect 505711 434094 505877 434110
rect 505911 434094 505978 434128
rect 506012 434094 506181 434128
rect 505711 434088 506181 434094
rect 505711 434054 506128 434088
rect 506162 434054 506181 434088
rect 505711 434020 505730 434054
rect 505764 434038 506181 434054
rect 505764 434020 505877 434038
rect 505711 434004 505877 434020
rect 505911 434004 505978 434038
rect 506012 434004 506181 434038
rect 505711 433998 506181 434004
rect 505711 433964 506128 433998
rect 506162 433964 506181 433998
rect 505711 433930 505730 433964
rect 505764 433948 506181 433964
rect 505764 433930 505877 433948
rect 505711 433914 505877 433930
rect 505911 433914 505978 433948
rect 506012 433914 506181 433948
rect 505711 433908 506181 433914
rect 505711 433874 506128 433908
rect 506162 433874 506181 433908
rect 505711 433840 505730 433874
rect 505764 433858 506181 433874
rect 505764 433840 505877 433858
rect 505711 433824 505877 433840
rect 505911 433824 505978 433858
rect 506012 433824 506181 433858
rect 505711 433818 506181 433824
rect 505711 433784 506128 433818
rect 506162 433784 506181 433818
rect 505711 433750 505730 433784
rect 505764 433768 506181 433784
rect 505764 433750 505877 433768
rect 505711 433734 505877 433750
rect 505911 433734 505978 433768
rect 506012 433734 506181 433768
rect 505711 433728 506181 433734
rect 505711 433694 506128 433728
rect 506162 433694 506181 433728
rect 505711 433660 505730 433694
rect 505764 433678 506181 433694
rect 505764 433660 505877 433678
rect 505711 433644 505877 433660
rect 505911 433644 505978 433678
rect 506012 433644 506181 433678
rect 505711 433638 506181 433644
rect 504423 433570 504442 433604
rect 504476 433588 504893 433604
rect 504476 433570 504589 433588
rect 504423 433565 504589 433570
rect 503436 433554 504589 433565
rect 504623 433554 504690 433588
rect 504724 433565 504893 433588
rect 505711 433604 506128 433638
rect 506162 433604 506181 433638
rect 506243 434260 506937 434321
rect 506243 434226 506304 434260
rect 506338 434248 506394 434260
rect 506428 434248 506484 434260
rect 506518 434248 506574 434260
rect 506350 434226 506394 434248
rect 506450 434226 506484 434248
rect 506550 434226 506574 434248
rect 506608 434248 506664 434260
rect 506608 434226 506616 434248
rect 506243 434214 506316 434226
rect 506350 434214 506416 434226
rect 506450 434214 506516 434226
rect 506550 434214 506616 434226
rect 506650 434226 506664 434248
rect 506698 434248 506754 434260
rect 506698 434226 506716 434248
rect 506650 434214 506716 434226
rect 506750 434226 506754 434248
rect 506788 434248 506844 434260
rect 506788 434226 506816 434248
rect 506878 434226 506937 434260
rect 506750 434214 506816 434226
rect 506850 434214 506937 434226
rect 506243 434170 506937 434214
rect 506243 434136 506304 434170
rect 506338 434148 506394 434170
rect 506428 434148 506484 434170
rect 506518 434148 506574 434170
rect 506350 434136 506394 434148
rect 506450 434136 506484 434148
rect 506550 434136 506574 434148
rect 506608 434148 506664 434170
rect 506608 434136 506616 434148
rect 506243 434114 506316 434136
rect 506350 434114 506416 434136
rect 506450 434114 506516 434136
rect 506550 434114 506616 434136
rect 506650 434136 506664 434148
rect 506698 434148 506754 434170
rect 506698 434136 506716 434148
rect 506650 434114 506716 434136
rect 506750 434136 506754 434148
rect 506788 434148 506844 434170
rect 506788 434136 506816 434148
rect 506878 434136 506937 434170
rect 506750 434114 506816 434136
rect 506850 434114 506937 434136
rect 506243 434080 506937 434114
rect 506243 434046 506304 434080
rect 506338 434048 506394 434080
rect 506428 434048 506484 434080
rect 506518 434048 506574 434080
rect 506350 434046 506394 434048
rect 506450 434046 506484 434048
rect 506550 434046 506574 434048
rect 506608 434048 506664 434080
rect 506608 434046 506616 434048
rect 506243 434014 506316 434046
rect 506350 434014 506416 434046
rect 506450 434014 506516 434046
rect 506550 434014 506616 434046
rect 506650 434046 506664 434048
rect 506698 434048 506754 434080
rect 506698 434046 506716 434048
rect 506650 434014 506716 434046
rect 506750 434046 506754 434048
rect 506788 434048 506844 434080
rect 506788 434046 506816 434048
rect 506878 434046 506937 434080
rect 506750 434014 506816 434046
rect 506850 434014 506937 434046
rect 506243 433990 506937 434014
rect 506243 433956 506304 433990
rect 506338 433956 506394 433990
rect 506428 433956 506484 433990
rect 506518 433956 506574 433990
rect 506608 433956 506664 433990
rect 506698 433956 506754 433990
rect 506788 433956 506844 433990
rect 506878 433956 506937 433990
rect 506243 433948 506937 433956
rect 506243 433914 506316 433948
rect 506350 433914 506416 433948
rect 506450 433914 506516 433948
rect 506550 433914 506616 433948
rect 506650 433914 506716 433948
rect 506750 433914 506816 433948
rect 506850 433914 506937 433948
rect 506243 433900 506937 433914
rect 506243 433866 506304 433900
rect 506338 433866 506394 433900
rect 506428 433866 506484 433900
rect 506518 433866 506574 433900
rect 506608 433866 506664 433900
rect 506698 433866 506754 433900
rect 506788 433866 506844 433900
rect 506878 433866 506937 433900
rect 506243 433848 506937 433866
rect 506243 433814 506316 433848
rect 506350 433814 506416 433848
rect 506450 433814 506516 433848
rect 506550 433814 506616 433848
rect 506650 433814 506716 433848
rect 506750 433814 506816 433848
rect 506850 433814 506937 433848
rect 506243 433810 506937 433814
rect 506243 433776 506304 433810
rect 506338 433776 506394 433810
rect 506428 433776 506484 433810
rect 506518 433776 506574 433810
rect 506608 433776 506664 433810
rect 506698 433776 506754 433810
rect 506788 433776 506844 433810
rect 506878 433776 506937 433810
rect 506243 433748 506937 433776
rect 506243 433720 506316 433748
rect 506350 433720 506416 433748
rect 506450 433720 506516 433748
rect 506550 433720 506616 433748
rect 506243 433686 506304 433720
rect 506350 433714 506394 433720
rect 506450 433714 506484 433720
rect 506550 433714 506574 433720
rect 506338 433686 506394 433714
rect 506428 433686 506484 433714
rect 506518 433686 506574 433714
rect 506608 433714 506616 433720
rect 506650 433720 506716 433748
rect 506650 433714 506664 433720
rect 506608 433686 506664 433714
rect 506698 433714 506716 433720
rect 506750 433720 506816 433748
rect 506850 433720 506937 433748
rect 506750 433714 506754 433720
rect 506698 433686 506754 433714
rect 506788 433714 506816 433720
rect 506788 433686 506844 433714
rect 506878 433686 506937 433720
rect 506243 433627 506937 433686
rect 506999 434290 507018 434324
rect 507052 434308 507469 434324
rect 508287 434364 508453 434383
rect 508487 434364 508554 434398
rect 508588 434383 509741 434398
rect 508588 434364 508757 434383
rect 508287 434358 508757 434364
rect 508287 434324 508704 434358
rect 508738 434324 508757 434358
rect 507052 434290 507165 434308
rect 506999 434274 507165 434290
rect 507199 434274 507266 434308
rect 507300 434274 507469 434308
rect 506999 434268 507469 434274
rect 506999 434234 507416 434268
rect 507450 434234 507469 434268
rect 506999 434200 507018 434234
rect 507052 434218 507469 434234
rect 507052 434200 507165 434218
rect 506999 434184 507165 434200
rect 507199 434184 507266 434218
rect 507300 434184 507469 434218
rect 506999 434178 507469 434184
rect 506999 434144 507416 434178
rect 507450 434144 507469 434178
rect 506999 434110 507018 434144
rect 507052 434128 507469 434144
rect 507052 434110 507165 434128
rect 506999 434094 507165 434110
rect 507199 434094 507266 434128
rect 507300 434094 507469 434128
rect 506999 434088 507469 434094
rect 506999 434054 507416 434088
rect 507450 434054 507469 434088
rect 506999 434020 507018 434054
rect 507052 434038 507469 434054
rect 507052 434020 507165 434038
rect 506999 434004 507165 434020
rect 507199 434004 507266 434038
rect 507300 434004 507469 434038
rect 506999 433998 507469 434004
rect 506999 433964 507416 433998
rect 507450 433964 507469 433998
rect 506999 433930 507018 433964
rect 507052 433948 507469 433964
rect 507052 433930 507165 433948
rect 506999 433914 507165 433930
rect 507199 433914 507266 433948
rect 507300 433914 507469 433948
rect 506999 433908 507469 433914
rect 506999 433874 507416 433908
rect 507450 433874 507469 433908
rect 506999 433840 507018 433874
rect 507052 433858 507469 433874
rect 507052 433840 507165 433858
rect 506999 433824 507165 433840
rect 507199 433824 507266 433858
rect 507300 433824 507469 433858
rect 506999 433818 507469 433824
rect 506999 433784 507416 433818
rect 507450 433784 507469 433818
rect 506999 433750 507018 433784
rect 507052 433768 507469 433784
rect 507052 433750 507165 433768
rect 506999 433734 507165 433750
rect 507199 433734 507266 433768
rect 507300 433734 507469 433768
rect 506999 433728 507469 433734
rect 506999 433694 507416 433728
rect 507450 433694 507469 433728
rect 506999 433660 507018 433694
rect 507052 433678 507469 433694
rect 507052 433660 507165 433678
rect 506999 433644 507165 433660
rect 507199 433644 507266 433678
rect 507300 433644 507469 433678
rect 506999 433638 507469 433644
rect 505711 433570 505730 433604
rect 505764 433588 506181 433604
rect 505764 433570 505877 433588
rect 505711 433565 505877 433570
rect 504724 433554 505877 433565
rect 505911 433554 505978 433588
rect 506012 433565 506181 433588
rect 506999 433604 507416 433638
rect 507450 433604 507469 433638
rect 507531 434260 508225 434321
rect 507531 434226 507592 434260
rect 507626 434248 507682 434260
rect 507716 434248 507772 434260
rect 507806 434248 507862 434260
rect 507638 434226 507682 434248
rect 507738 434226 507772 434248
rect 507838 434226 507862 434248
rect 507896 434248 507952 434260
rect 507896 434226 507904 434248
rect 507531 434214 507604 434226
rect 507638 434214 507704 434226
rect 507738 434214 507804 434226
rect 507838 434214 507904 434226
rect 507938 434226 507952 434248
rect 507986 434248 508042 434260
rect 507986 434226 508004 434248
rect 507938 434214 508004 434226
rect 508038 434226 508042 434248
rect 508076 434248 508132 434260
rect 508076 434226 508104 434248
rect 508166 434226 508225 434260
rect 508038 434214 508104 434226
rect 508138 434214 508225 434226
rect 507531 434170 508225 434214
rect 507531 434136 507592 434170
rect 507626 434148 507682 434170
rect 507716 434148 507772 434170
rect 507806 434148 507862 434170
rect 507638 434136 507682 434148
rect 507738 434136 507772 434148
rect 507838 434136 507862 434148
rect 507896 434148 507952 434170
rect 507896 434136 507904 434148
rect 507531 434114 507604 434136
rect 507638 434114 507704 434136
rect 507738 434114 507804 434136
rect 507838 434114 507904 434136
rect 507938 434136 507952 434148
rect 507986 434148 508042 434170
rect 507986 434136 508004 434148
rect 507938 434114 508004 434136
rect 508038 434136 508042 434148
rect 508076 434148 508132 434170
rect 508076 434136 508104 434148
rect 508166 434136 508225 434170
rect 508038 434114 508104 434136
rect 508138 434114 508225 434136
rect 507531 434080 508225 434114
rect 507531 434046 507592 434080
rect 507626 434048 507682 434080
rect 507716 434048 507772 434080
rect 507806 434048 507862 434080
rect 507638 434046 507682 434048
rect 507738 434046 507772 434048
rect 507838 434046 507862 434048
rect 507896 434048 507952 434080
rect 507896 434046 507904 434048
rect 507531 434014 507604 434046
rect 507638 434014 507704 434046
rect 507738 434014 507804 434046
rect 507838 434014 507904 434046
rect 507938 434046 507952 434048
rect 507986 434048 508042 434080
rect 507986 434046 508004 434048
rect 507938 434014 508004 434046
rect 508038 434046 508042 434048
rect 508076 434048 508132 434080
rect 508076 434046 508104 434048
rect 508166 434046 508225 434080
rect 508038 434014 508104 434046
rect 508138 434014 508225 434046
rect 507531 433990 508225 434014
rect 507531 433956 507592 433990
rect 507626 433956 507682 433990
rect 507716 433956 507772 433990
rect 507806 433956 507862 433990
rect 507896 433956 507952 433990
rect 507986 433956 508042 433990
rect 508076 433956 508132 433990
rect 508166 433956 508225 433990
rect 507531 433948 508225 433956
rect 507531 433914 507604 433948
rect 507638 433914 507704 433948
rect 507738 433914 507804 433948
rect 507838 433914 507904 433948
rect 507938 433914 508004 433948
rect 508038 433914 508104 433948
rect 508138 433914 508225 433948
rect 507531 433900 508225 433914
rect 507531 433866 507592 433900
rect 507626 433866 507682 433900
rect 507716 433866 507772 433900
rect 507806 433866 507862 433900
rect 507896 433866 507952 433900
rect 507986 433866 508042 433900
rect 508076 433866 508132 433900
rect 508166 433866 508225 433900
rect 507531 433848 508225 433866
rect 507531 433814 507604 433848
rect 507638 433814 507704 433848
rect 507738 433814 507804 433848
rect 507838 433814 507904 433848
rect 507938 433814 508004 433848
rect 508038 433814 508104 433848
rect 508138 433814 508225 433848
rect 507531 433810 508225 433814
rect 507531 433776 507592 433810
rect 507626 433776 507682 433810
rect 507716 433776 507772 433810
rect 507806 433776 507862 433810
rect 507896 433776 507952 433810
rect 507986 433776 508042 433810
rect 508076 433776 508132 433810
rect 508166 433776 508225 433810
rect 507531 433748 508225 433776
rect 507531 433720 507604 433748
rect 507638 433720 507704 433748
rect 507738 433720 507804 433748
rect 507838 433720 507904 433748
rect 507531 433686 507592 433720
rect 507638 433714 507682 433720
rect 507738 433714 507772 433720
rect 507838 433714 507862 433720
rect 507626 433686 507682 433714
rect 507716 433686 507772 433714
rect 507806 433686 507862 433714
rect 507896 433714 507904 433720
rect 507938 433720 508004 433748
rect 507938 433714 507952 433720
rect 507896 433686 507952 433714
rect 507986 433714 508004 433720
rect 508038 433720 508104 433748
rect 508138 433720 508225 433748
rect 508038 433714 508042 433720
rect 507986 433686 508042 433714
rect 508076 433714 508104 433720
rect 508076 433686 508132 433714
rect 508166 433686 508225 433720
rect 507531 433627 508225 433686
rect 508287 434290 508306 434324
rect 508340 434308 508757 434324
rect 509575 434364 509741 434383
rect 509775 434364 509842 434398
rect 509876 434383 511029 434398
rect 509876 434364 510045 434383
rect 509575 434358 510045 434364
rect 509575 434324 509992 434358
rect 510026 434324 510045 434358
rect 508340 434290 508453 434308
rect 508287 434274 508453 434290
rect 508487 434274 508554 434308
rect 508588 434274 508757 434308
rect 508287 434268 508757 434274
rect 508287 434234 508704 434268
rect 508738 434234 508757 434268
rect 508287 434200 508306 434234
rect 508340 434218 508757 434234
rect 508340 434200 508453 434218
rect 508287 434184 508453 434200
rect 508487 434184 508554 434218
rect 508588 434184 508757 434218
rect 508287 434178 508757 434184
rect 508287 434144 508704 434178
rect 508738 434144 508757 434178
rect 508287 434110 508306 434144
rect 508340 434128 508757 434144
rect 508340 434110 508453 434128
rect 508287 434094 508453 434110
rect 508487 434094 508554 434128
rect 508588 434094 508757 434128
rect 508287 434088 508757 434094
rect 508287 434054 508704 434088
rect 508738 434054 508757 434088
rect 508287 434020 508306 434054
rect 508340 434038 508757 434054
rect 508340 434020 508453 434038
rect 508287 434004 508453 434020
rect 508487 434004 508554 434038
rect 508588 434004 508757 434038
rect 508287 433998 508757 434004
rect 508287 433964 508704 433998
rect 508738 433964 508757 433998
rect 508287 433930 508306 433964
rect 508340 433948 508757 433964
rect 508340 433930 508453 433948
rect 508287 433914 508453 433930
rect 508487 433914 508554 433948
rect 508588 433914 508757 433948
rect 508287 433908 508757 433914
rect 508287 433874 508704 433908
rect 508738 433874 508757 433908
rect 508287 433840 508306 433874
rect 508340 433858 508757 433874
rect 508340 433840 508453 433858
rect 508287 433824 508453 433840
rect 508487 433824 508554 433858
rect 508588 433824 508757 433858
rect 508287 433818 508757 433824
rect 508287 433784 508704 433818
rect 508738 433784 508757 433818
rect 508287 433750 508306 433784
rect 508340 433768 508757 433784
rect 508340 433750 508453 433768
rect 508287 433734 508453 433750
rect 508487 433734 508554 433768
rect 508588 433734 508757 433768
rect 508287 433728 508757 433734
rect 508287 433694 508704 433728
rect 508738 433694 508757 433728
rect 508287 433660 508306 433694
rect 508340 433678 508757 433694
rect 508340 433660 508453 433678
rect 508287 433644 508453 433660
rect 508487 433644 508554 433678
rect 508588 433644 508757 433678
rect 508287 433638 508757 433644
rect 506999 433570 507018 433604
rect 507052 433588 507469 433604
rect 507052 433570 507165 433588
rect 506999 433565 507165 433570
rect 506012 433554 507165 433565
rect 507199 433554 507266 433588
rect 507300 433565 507469 433588
rect 508287 433604 508704 433638
rect 508738 433604 508757 433638
rect 508819 434260 509513 434321
rect 508819 434226 508880 434260
rect 508914 434248 508970 434260
rect 509004 434248 509060 434260
rect 509094 434248 509150 434260
rect 508926 434226 508970 434248
rect 509026 434226 509060 434248
rect 509126 434226 509150 434248
rect 509184 434248 509240 434260
rect 509184 434226 509192 434248
rect 508819 434214 508892 434226
rect 508926 434214 508992 434226
rect 509026 434214 509092 434226
rect 509126 434214 509192 434226
rect 509226 434226 509240 434248
rect 509274 434248 509330 434260
rect 509274 434226 509292 434248
rect 509226 434214 509292 434226
rect 509326 434226 509330 434248
rect 509364 434248 509420 434260
rect 509364 434226 509392 434248
rect 509454 434226 509513 434260
rect 509326 434214 509392 434226
rect 509426 434214 509513 434226
rect 508819 434170 509513 434214
rect 508819 434136 508880 434170
rect 508914 434148 508970 434170
rect 509004 434148 509060 434170
rect 509094 434148 509150 434170
rect 508926 434136 508970 434148
rect 509026 434136 509060 434148
rect 509126 434136 509150 434148
rect 509184 434148 509240 434170
rect 509184 434136 509192 434148
rect 508819 434114 508892 434136
rect 508926 434114 508992 434136
rect 509026 434114 509092 434136
rect 509126 434114 509192 434136
rect 509226 434136 509240 434148
rect 509274 434148 509330 434170
rect 509274 434136 509292 434148
rect 509226 434114 509292 434136
rect 509326 434136 509330 434148
rect 509364 434148 509420 434170
rect 509364 434136 509392 434148
rect 509454 434136 509513 434170
rect 509326 434114 509392 434136
rect 509426 434114 509513 434136
rect 508819 434080 509513 434114
rect 508819 434046 508880 434080
rect 508914 434048 508970 434080
rect 509004 434048 509060 434080
rect 509094 434048 509150 434080
rect 508926 434046 508970 434048
rect 509026 434046 509060 434048
rect 509126 434046 509150 434048
rect 509184 434048 509240 434080
rect 509184 434046 509192 434048
rect 508819 434014 508892 434046
rect 508926 434014 508992 434046
rect 509026 434014 509092 434046
rect 509126 434014 509192 434046
rect 509226 434046 509240 434048
rect 509274 434048 509330 434080
rect 509274 434046 509292 434048
rect 509226 434014 509292 434046
rect 509326 434046 509330 434048
rect 509364 434048 509420 434080
rect 509364 434046 509392 434048
rect 509454 434046 509513 434080
rect 509326 434014 509392 434046
rect 509426 434014 509513 434046
rect 508819 433990 509513 434014
rect 508819 433956 508880 433990
rect 508914 433956 508970 433990
rect 509004 433956 509060 433990
rect 509094 433956 509150 433990
rect 509184 433956 509240 433990
rect 509274 433956 509330 433990
rect 509364 433956 509420 433990
rect 509454 433956 509513 433990
rect 508819 433948 509513 433956
rect 508819 433914 508892 433948
rect 508926 433914 508992 433948
rect 509026 433914 509092 433948
rect 509126 433914 509192 433948
rect 509226 433914 509292 433948
rect 509326 433914 509392 433948
rect 509426 433914 509513 433948
rect 508819 433900 509513 433914
rect 508819 433866 508880 433900
rect 508914 433866 508970 433900
rect 509004 433866 509060 433900
rect 509094 433866 509150 433900
rect 509184 433866 509240 433900
rect 509274 433866 509330 433900
rect 509364 433866 509420 433900
rect 509454 433866 509513 433900
rect 508819 433848 509513 433866
rect 508819 433814 508892 433848
rect 508926 433814 508992 433848
rect 509026 433814 509092 433848
rect 509126 433814 509192 433848
rect 509226 433814 509292 433848
rect 509326 433814 509392 433848
rect 509426 433814 509513 433848
rect 508819 433810 509513 433814
rect 508819 433776 508880 433810
rect 508914 433776 508970 433810
rect 509004 433776 509060 433810
rect 509094 433776 509150 433810
rect 509184 433776 509240 433810
rect 509274 433776 509330 433810
rect 509364 433776 509420 433810
rect 509454 433776 509513 433810
rect 508819 433748 509513 433776
rect 508819 433720 508892 433748
rect 508926 433720 508992 433748
rect 509026 433720 509092 433748
rect 509126 433720 509192 433748
rect 508819 433686 508880 433720
rect 508926 433714 508970 433720
rect 509026 433714 509060 433720
rect 509126 433714 509150 433720
rect 508914 433686 508970 433714
rect 509004 433686 509060 433714
rect 509094 433686 509150 433714
rect 509184 433714 509192 433720
rect 509226 433720 509292 433748
rect 509226 433714 509240 433720
rect 509184 433686 509240 433714
rect 509274 433714 509292 433720
rect 509326 433720 509392 433748
rect 509426 433720 509513 433748
rect 509326 433714 509330 433720
rect 509274 433686 509330 433714
rect 509364 433714 509392 433720
rect 509364 433686 509420 433714
rect 509454 433686 509513 433720
rect 508819 433627 509513 433686
rect 509575 434290 509594 434324
rect 509628 434308 510045 434324
rect 510863 434364 511029 434383
rect 511063 434364 511130 434398
rect 511164 434383 512317 434398
rect 511164 434364 511333 434383
rect 510863 434358 511333 434364
rect 510863 434324 511280 434358
rect 511314 434324 511333 434358
rect 509628 434290 509741 434308
rect 509575 434274 509741 434290
rect 509775 434274 509842 434308
rect 509876 434274 510045 434308
rect 509575 434268 510045 434274
rect 509575 434234 509992 434268
rect 510026 434234 510045 434268
rect 509575 434200 509594 434234
rect 509628 434218 510045 434234
rect 509628 434200 509741 434218
rect 509575 434184 509741 434200
rect 509775 434184 509842 434218
rect 509876 434184 510045 434218
rect 509575 434178 510045 434184
rect 509575 434144 509992 434178
rect 510026 434144 510045 434178
rect 509575 434110 509594 434144
rect 509628 434128 510045 434144
rect 509628 434110 509741 434128
rect 509575 434094 509741 434110
rect 509775 434094 509842 434128
rect 509876 434094 510045 434128
rect 509575 434088 510045 434094
rect 509575 434054 509992 434088
rect 510026 434054 510045 434088
rect 509575 434020 509594 434054
rect 509628 434038 510045 434054
rect 509628 434020 509741 434038
rect 509575 434004 509741 434020
rect 509775 434004 509842 434038
rect 509876 434004 510045 434038
rect 509575 433998 510045 434004
rect 509575 433964 509992 433998
rect 510026 433964 510045 433998
rect 509575 433930 509594 433964
rect 509628 433948 510045 433964
rect 509628 433930 509741 433948
rect 509575 433914 509741 433930
rect 509775 433914 509842 433948
rect 509876 433914 510045 433948
rect 509575 433908 510045 433914
rect 509575 433874 509992 433908
rect 510026 433874 510045 433908
rect 509575 433840 509594 433874
rect 509628 433858 510045 433874
rect 509628 433840 509741 433858
rect 509575 433824 509741 433840
rect 509775 433824 509842 433858
rect 509876 433824 510045 433858
rect 509575 433818 510045 433824
rect 509575 433784 509992 433818
rect 510026 433784 510045 433818
rect 509575 433750 509594 433784
rect 509628 433768 510045 433784
rect 509628 433750 509741 433768
rect 509575 433734 509741 433750
rect 509775 433734 509842 433768
rect 509876 433734 510045 433768
rect 509575 433728 510045 433734
rect 509575 433694 509992 433728
rect 510026 433694 510045 433728
rect 509575 433660 509594 433694
rect 509628 433678 510045 433694
rect 509628 433660 509741 433678
rect 509575 433644 509741 433660
rect 509775 433644 509842 433678
rect 509876 433644 510045 433678
rect 509575 433638 510045 433644
rect 508287 433570 508306 433604
rect 508340 433588 508757 433604
rect 508340 433570 508453 433588
rect 508287 433565 508453 433570
rect 507300 433554 508453 433565
rect 508487 433554 508554 433588
rect 508588 433565 508757 433588
rect 509575 433604 509992 433638
rect 510026 433604 510045 433638
rect 510107 434260 510801 434321
rect 510107 434226 510168 434260
rect 510202 434248 510258 434260
rect 510292 434248 510348 434260
rect 510382 434248 510438 434260
rect 510214 434226 510258 434248
rect 510314 434226 510348 434248
rect 510414 434226 510438 434248
rect 510472 434248 510528 434260
rect 510472 434226 510480 434248
rect 510107 434214 510180 434226
rect 510214 434214 510280 434226
rect 510314 434214 510380 434226
rect 510414 434214 510480 434226
rect 510514 434226 510528 434248
rect 510562 434248 510618 434260
rect 510562 434226 510580 434248
rect 510514 434214 510580 434226
rect 510614 434226 510618 434248
rect 510652 434248 510708 434260
rect 510652 434226 510680 434248
rect 510742 434226 510801 434260
rect 510614 434214 510680 434226
rect 510714 434214 510801 434226
rect 510107 434170 510801 434214
rect 510107 434136 510168 434170
rect 510202 434148 510258 434170
rect 510292 434148 510348 434170
rect 510382 434148 510438 434170
rect 510214 434136 510258 434148
rect 510314 434136 510348 434148
rect 510414 434136 510438 434148
rect 510472 434148 510528 434170
rect 510472 434136 510480 434148
rect 510107 434114 510180 434136
rect 510214 434114 510280 434136
rect 510314 434114 510380 434136
rect 510414 434114 510480 434136
rect 510514 434136 510528 434148
rect 510562 434148 510618 434170
rect 510562 434136 510580 434148
rect 510514 434114 510580 434136
rect 510614 434136 510618 434148
rect 510652 434148 510708 434170
rect 510652 434136 510680 434148
rect 510742 434136 510801 434170
rect 510614 434114 510680 434136
rect 510714 434114 510801 434136
rect 510107 434080 510801 434114
rect 510107 434046 510168 434080
rect 510202 434048 510258 434080
rect 510292 434048 510348 434080
rect 510382 434048 510438 434080
rect 510214 434046 510258 434048
rect 510314 434046 510348 434048
rect 510414 434046 510438 434048
rect 510472 434048 510528 434080
rect 510472 434046 510480 434048
rect 510107 434014 510180 434046
rect 510214 434014 510280 434046
rect 510314 434014 510380 434046
rect 510414 434014 510480 434046
rect 510514 434046 510528 434048
rect 510562 434048 510618 434080
rect 510562 434046 510580 434048
rect 510514 434014 510580 434046
rect 510614 434046 510618 434048
rect 510652 434048 510708 434080
rect 510652 434046 510680 434048
rect 510742 434046 510801 434080
rect 510614 434014 510680 434046
rect 510714 434014 510801 434046
rect 510107 433990 510801 434014
rect 510107 433956 510168 433990
rect 510202 433956 510258 433990
rect 510292 433956 510348 433990
rect 510382 433956 510438 433990
rect 510472 433956 510528 433990
rect 510562 433956 510618 433990
rect 510652 433956 510708 433990
rect 510742 433956 510801 433990
rect 510107 433948 510801 433956
rect 510107 433914 510180 433948
rect 510214 433914 510280 433948
rect 510314 433914 510380 433948
rect 510414 433914 510480 433948
rect 510514 433914 510580 433948
rect 510614 433914 510680 433948
rect 510714 433914 510801 433948
rect 510107 433900 510801 433914
rect 510107 433866 510168 433900
rect 510202 433866 510258 433900
rect 510292 433866 510348 433900
rect 510382 433866 510438 433900
rect 510472 433866 510528 433900
rect 510562 433866 510618 433900
rect 510652 433866 510708 433900
rect 510742 433866 510801 433900
rect 510107 433848 510801 433866
rect 510107 433814 510180 433848
rect 510214 433814 510280 433848
rect 510314 433814 510380 433848
rect 510414 433814 510480 433848
rect 510514 433814 510580 433848
rect 510614 433814 510680 433848
rect 510714 433814 510801 433848
rect 510107 433810 510801 433814
rect 510107 433776 510168 433810
rect 510202 433776 510258 433810
rect 510292 433776 510348 433810
rect 510382 433776 510438 433810
rect 510472 433776 510528 433810
rect 510562 433776 510618 433810
rect 510652 433776 510708 433810
rect 510742 433776 510801 433810
rect 510107 433748 510801 433776
rect 510107 433720 510180 433748
rect 510214 433720 510280 433748
rect 510314 433720 510380 433748
rect 510414 433720 510480 433748
rect 510107 433686 510168 433720
rect 510214 433714 510258 433720
rect 510314 433714 510348 433720
rect 510414 433714 510438 433720
rect 510202 433686 510258 433714
rect 510292 433686 510348 433714
rect 510382 433686 510438 433714
rect 510472 433714 510480 433720
rect 510514 433720 510580 433748
rect 510514 433714 510528 433720
rect 510472 433686 510528 433714
rect 510562 433714 510580 433720
rect 510614 433720 510680 433748
rect 510714 433720 510801 433748
rect 510614 433714 510618 433720
rect 510562 433686 510618 433714
rect 510652 433714 510680 433720
rect 510652 433686 510708 433714
rect 510742 433686 510801 433720
rect 510107 433627 510801 433686
rect 510863 434290 510882 434324
rect 510916 434308 511333 434324
rect 512151 434364 512317 434383
rect 512351 434364 512418 434398
rect 512452 434383 513605 434398
rect 512452 434364 512621 434383
rect 512151 434358 512621 434364
rect 512151 434324 512568 434358
rect 512602 434324 512621 434358
rect 510916 434290 511029 434308
rect 510863 434274 511029 434290
rect 511063 434274 511130 434308
rect 511164 434274 511333 434308
rect 510863 434268 511333 434274
rect 510863 434234 511280 434268
rect 511314 434234 511333 434268
rect 510863 434200 510882 434234
rect 510916 434218 511333 434234
rect 510916 434200 511029 434218
rect 510863 434184 511029 434200
rect 511063 434184 511130 434218
rect 511164 434184 511333 434218
rect 510863 434178 511333 434184
rect 510863 434144 511280 434178
rect 511314 434144 511333 434178
rect 510863 434110 510882 434144
rect 510916 434128 511333 434144
rect 510916 434110 511029 434128
rect 510863 434094 511029 434110
rect 511063 434094 511130 434128
rect 511164 434094 511333 434128
rect 510863 434088 511333 434094
rect 510863 434054 511280 434088
rect 511314 434054 511333 434088
rect 510863 434020 510882 434054
rect 510916 434038 511333 434054
rect 510916 434020 511029 434038
rect 510863 434004 511029 434020
rect 511063 434004 511130 434038
rect 511164 434004 511333 434038
rect 510863 433998 511333 434004
rect 510863 433964 511280 433998
rect 511314 433964 511333 433998
rect 510863 433930 510882 433964
rect 510916 433948 511333 433964
rect 510916 433930 511029 433948
rect 510863 433914 511029 433930
rect 511063 433914 511130 433948
rect 511164 433914 511333 433948
rect 510863 433908 511333 433914
rect 510863 433874 511280 433908
rect 511314 433874 511333 433908
rect 510863 433840 510882 433874
rect 510916 433858 511333 433874
rect 510916 433840 511029 433858
rect 510863 433824 511029 433840
rect 511063 433824 511130 433858
rect 511164 433824 511333 433858
rect 510863 433818 511333 433824
rect 510863 433784 511280 433818
rect 511314 433784 511333 433818
rect 510863 433750 510882 433784
rect 510916 433768 511333 433784
rect 510916 433750 511029 433768
rect 510863 433734 511029 433750
rect 511063 433734 511130 433768
rect 511164 433734 511333 433768
rect 510863 433728 511333 433734
rect 510863 433694 511280 433728
rect 511314 433694 511333 433728
rect 510863 433660 510882 433694
rect 510916 433678 511333 433694
rect 510916 433660 511029 433678
rect 510863 433644 511029 433660
rect 511063 433644 511130 433678
rect 511164 433644 511333 433678
rect 510863 433638 511333 433644
rect 509575 433570 509594 433604
rect 509628 433588 510045 433604
rect 509628 433570 509741 433588
rect 509575 433565 509741 433570
rect 508588 433554 509741 433565
rect 509775 433554 509842 433588
rect 509876 433565 510045 433588
rect 510863 433604 511280 433638
rect 511314 433604 511333 433638
rect 511395 434260 512089 434321
rect 511395 434226 511456 434260
rect 511490 434248 511546 434260
rect 511580 434248 511636 434260
rect 511670 434248 511726 434260
rect 511502 434226 511546 434248
rect 511602 434226 511636 434248
rect 511702 434226 511726 434248
rect 511760 434248 511816 434260
rect 511760 434226 511768 434248
rect 511395 434214 511468 434226
rect 511502 434214 511568 434226
rect 511602 434214 511668 434226
rect 511702 434214 511768 434226
rect 511802 434226 511816 434248
rect 511850 434248 511906 434260
rect 511850 434226 511868 434248
rect 511802 434214 511868 434226
rect 511902 434226 511906 434248
rect 511940 434248 511996 434260
rect 511940 434226 511968 434248
rect 512030 434226 512089 434260
rect 511902 434214 511968 434226
rect 512002 434214 512089 434226
rect 511395 434170 512089 434214
rect 511395 434136 511456 434170
rect 511490 434148 511546 434170
rect 511580 434148 511636 434170
rect 511670 434148 511726 434170
rect 511502 434136 511546 434148
rect 511602 434136 511636 434148
rect 511702 434136 511726 434148
rect 511760 434148 511816 434170
rect 511760 434136 511768 434148
rect 511395 434114 511468 434136
rect 511502 434114 511568 434136
rect 511602 434114 511668 434136
rect 511702 434114 511768 434136
rect 511802 434136 511816 434148
rect 511850 434148 511906 434170
rect 511850 434136 511868 434148
rect 511802 434114 511868 434136
rect 511902 434136 511906 434148
rect 511940 434148 511996 434170
rect 511940 434136 511968 434148
rect 512030 434136 512089 434170
rect 511902 434114 511968 434136
rect 512002 434114 512089 434136
rect 511395 434080 512089 434114
rect 511395 434046 511456 434080
rect 511490 434048 511546 434080
rect 511580 434048 511636 434080
rect 511670 434048 511726 434080
rect 511502 434046 511546 434048
rect 511602 434046 511636 434048
rect 511702 434046 511726 434048
rect 511760 434048 511816 434080
rect 511760 434046 511768 434048
rect 511395 434014 511468 434046
rect 511502 434014 511568 434046
rect 511602 434014 511668 434046
rect 511702 434014 511768 434046
rect 511802 434046 511816 434048
rect 511850 434048 511906 434080
rect 511850 434046 511868 434048
rect 511802 434014 511868 434046
rect 511902 434046 511906 434048
rect 511940 434048 511996 434080
rect 511940 434046 511968 434048
rect 512030 434046 512089 434080
rect 511902 434014 511968 434046
rect 512002 434014 512089 434046
rect 511395 433990 512089 434014
rect 511395 433956 511456 433990
rect 511490 433956 511546 433990
rect 511580 433956 511636 433990
rect 511670 433956 511726 433990
rect 511760 433956 511816 433990
rect 511850 433956 511906 433990
rect 511940 433956 511996 433990
rect 512030 433956 512089 433990
rect 511395 433948 512089 433956
rect 511395 433914 511468 433948
rect 511502 433914 511568 433948
rect 511602 433914 511668 433948
rect 511702 433914 511768 433948
rect 511802 433914 511868 433948
rect 511902 433914 511968 433948
rect 512002 433914 512089 433948
rect 511395 433900 512089 433914
rect 511395 433866 511456 433900
rect 511490 433866 511546 433900
rect 511580 433866 511636 433900
rect 511670 433866 511726 433900
rect 511760 433866 511816 433900
rect 511850 433866 511906 433900
rect 511940 433866 511996 433900
rect 512030 433866 512089 433900
rect 511395 433848 512089 433866
rect 511395 433814 511468 433848
rect 511502 433814 511568 433848
rect 511602 433814 511668 433848
rect 511702 433814 511768 433848
rect 511802 433814 511868 433848
rect 511902 433814 511968 433848
rect 512002 433814 512089 433848
rect 511395 433810 512089 433814
rect 511395 433776 511456 433810
rect 511490 433776 511546 433810
rect 511580 433776 511636 433810
rect 511670 433776 511726 433810
rect 511760 433776 511816 433810
rect 511850 433776 511906 433810
rect 511940 433776 511996 433810
rect 512030 433776 512089 433810
rect 511395 433748 512089 433776
rect 511395 433720 511468 433748
rect 511502 433720 511568 433748
rect 511602 433720 511668 433748
rect 511702 433720 511768 433748
rect 511395 433686 511456 433720
rect 511502 433714 511546 433720
rect 511602 433714 511636 433720
rect 511702 433714 511726 433720
rect 511490 433686 511546 433714
rect 511580 433686 511636 433714
rect 511670 433686 511726 433714
rect 511760 433714 511768 433720
rect 511802 433720 511868 433748
rect 511802 433714 511816 433720
rect 511760 433686 511816 433714
rect 511850 433714 511868 433720
rect 511902 433720 511968 433748
rect 512002 433720 512089 433748
rect 511902 433714 511906 433720
rect 511850 433686 511906 433714
rect 511940 433714 511968 433720
rect 511940 433686 511996 433714
rect 512030 433686 512089 433720
rect 511395 433627 512089 433686
rect 512151 434290 512170 434324
rect 512204 434308 512621 434324
rect 513439 434364 513605 434383
rect 513639 434364 513674 434398
rect 513439 434324 513674 434364
rect 512204 434290 512317 434308
rect 512151 434274 512317 434290
rect 512351 434274 512418 434308
rect 512452 434274 512621 434308
rect 512151 434268 512621 434274
rect 512151 434234 512568 434268
rect 512602 434234 512621 434268
rect 512151 434200 512170 434234
rect 512204 434218 512621 434234
rect 512204 434200 512317 434218
rect 512151 434184 512317 434200
rect 512351 434184 512418 434218
rect 512452 434184 512621 434218
rect 512151 434178 512621 434184
rect 512151 434144 512568 434178
rect 512602 434144 512621 434178
rect 512151 434110 512170 434144
rect 512204 434128 512621 434144
rect 512204 434110 512317 434128
rect 512151 434094 512317 434110
rect 512351 434094 512418 434128
rect 512452 434094 512621 434128
rect 512151 434088 512621 434094
rect 512151 434054 512568 434088
rect 512602 434054 512621 434088
rect 512151 434020 512170 434054
rect 512204 434038 512621 434054
rect 512204 434020 512317 434038
rect 512151 434004 512317 434020
rect 512351 434004 512418 434038
rect 512452 434004 512621 434038
rect 512151 433998 512621 434004
rect 512151 433964 512568 433998
rect 512602 433964 512621 433998
rect 512151 433930 512170 433964
rect 512204 433948 512621 433964
rect 512204 433930 512317 433948
rect 512151 433914 512317 433930
rect 512351 433914 512418 433948
rect 512452 433914 512621 433948
rect 512151 433908 512621 433914
rect 512151 433874 512568 433908
rect 512602 433874 512621 433908
rect 512151 433840 512170 433874
rect 512204 433858 512621 433874
rect 512204 433840 512317 433858
rect 512151 433824 512317 433840
rect 512351 433824 512418 433858
rect 512452 433824 512621 433858
rect 512151 433818 512621 433824
rect 512151 433784 512568 433818
rect 512602 433784 512621 433818
rect 512151 433750 512170 433784
rect 512204 433768 512621 433784
rect 512204 433750 512317 433768
rect 512151 433734 512317 433750
rect 512351 433734 512418 433768
rect 512452 433734 512621 433768
rect 512151 433728 512621 433734
rect 512151 433694 512568 433728
rect 512602 433694 512621 433728
rect 512151 433660 512170 433694
rect 512204 433678 512621 433694
rect 512204 433660 512317 433678
rect 512151 433644 512317 433660
rect 512351 433644 512418 433678
rect 512452 433644 512621 433678
rect 512151 433638 512621 433644
rect 510863 433570 510882 433604
rect 510916 433588 511333 433604
rect 510916 433570 511029 433588
rect 510863 433565 511029 433570
rect 509876 433554 511029 433565
rect 511063 433554 511130 433588
rect 511164 433565 511333 433588
rect 512151 433604 512568 433638
rect 512602 433604 512621 433638
rect 512683 434260 513377 434321
rect 512683 434226 512744 434260
rect 512778 434248 512834 434260
rect 512868 434248 512924 434260
rect 512958 434248 513014 434260
rect 512790 434226 512834 434248
rect 512890 434226 512924 434248
rect 512990 434226 513014 434248
rect 513048 434248 513104 434260
rect 513048 434226 513056 434248
rect 512683 434214 512756 434226
rect 512790 434214 512856 434226
rect 512890 434214 512956 434226
rect 512990 434214 513056 434226
rect 513090 434226 513104 434248
rect 513138 434248 513194 434260
rect 513138 434226 513156 434248
rect 513090 434214 513156 434226
rect 513190 434226 513194 434248
rect 513228 434248 513284 434260
rect 513228 434226 513256 434248
rect 513318 434226 513377 434260
rect 513190 434214 513256 434226
rect 513290 434214 513377 434226
rect 512683 434170 513377 434214
rect 512683 434136 512744 434170
rect 512778 434148 512834 434170
rect 512868 434148 512924 434170
rect 512958 434148 513014 434170
rect 512790 434136 512834 434148
rect 512890 434136 512924 434148
rect 512990 434136 513014 434148
rect 513048 434148 513104 434170
rect 513048 434136 513056 434148
rect 512683 434114 512756 434136
rect 512790 434114 512856 434136
rect 512890 434114 512956 434136
rect 512990 434114 513056 434136
rect 513090 434136 513104 434148
rect 513138 434148 513194 434170
rect 513138 434136 513156 434148
rect 513090 434114 513156 434136
rect 513190 434136 513194 434148
rect 513228 434148 513284 434170
rect 513228 434136 513256 434148
rect 513318 434136 513377 434170
rect 513190 434114 513256 434136
rect 513290 434114 513377 434136
rect 512683 434080 513377 434114
rect 512683 434046 512744 434080
rect 512778 434048 512834 434080
rect 512868 434048 512924 434080
rect 512958 434048 513014 434080
rect 512790 434046 512834 434048
rect 512890 434046 512924 434048
rect 512990 434046 513014 434048
rect 513048 434048 513104 434080
rect 513048 434046 513056 434048
rect 512683 434014 512756 434046
rect 512790 434014 512856 434046
rect 512890 434014 512956 434046
rect 512990 434014 513056 434046
rect 513090 434046 513104 434048
rect 513138 434048 513194 434080
rect 513138 434046 513156 434048
rect 513090 434014 513156 434046
rect 513190 434046 513194 434048
rect 513228 434048 513284 434080
rect 513228 434046 513256 434048
rect 513318 434046 513377 434080
rect 513190 434014 513256 434046
rect 513290 434014 513377 434046
rect 512683 433990 513377 434014
rect 512683 433956 512744 433990
rect 512778 433956 512834 433990
rect 512868 433956 512924 433990
rect 512958 433956 513014 433990
rect 513048 433956 513104 433990
rect 513138 433956 513194 433990
rect 513228 433956 513284 433990
rect 513318 433956 513377 433990
rect 512683 433948 513377 433956
rect 512683 433914 512756 433948
rect 512790 433914 512856 433948
rect 512890 433914 512956 433948
rect 512990 433914 513056 433948
rect 513090 433914 513156 433948
rect 513190 433914 513256 433948
rect 513290 433914 513377 433948
rect 512683 433900 513377 433914
rect 512683 433866 512744 433900
rect 512778 433866 512834 433900
rect 512868 433866 512924 433900
rect 512958 433866 513014 433900
rect 513048 433866 513104 433900
rect 513138 433866 513194 433900
rect 513228 433866 513284 433900
rect 513318 433866 513377 433900
rect 512683 433848 513377 433866
rect 512683 433814 512756 433848
rect 512790 433814 512856 433848
rect 512890 433814 512956 433848
rect 512990 433814 513056 433848
rect 513090 433814 513156 433848
rect 513190 433814 513256 433848
rect 513290 433814 513377 433848
rect 512683 433810 513377 433814
rect 512683 433776 512744 433810
rect 512778 433776 512834 433810
rect 512868 433776 512924 433810
rect 512958 433776 513014 433810
rect 513048 433776 513104 433810
rect 513138 433776 513194 433810
rect 513228 433776 513284 433810
rect 513318 433776 513377 433810
rect 512683 433748 513377 433776
rect 512683 433720 512756 433748
rect 512790 433720 512856 433748
rect 512890 433720 512956 433748
rect 512990 433720 513056 433748
rect 512683 433686 512744 433720
rect 512790 433714 512834 433720
rect 512890 433714 512924 433720
rect 512990 433714 513014 433720
rect 512778 433686 512834 433714
rect 512868 433686 512924 433714
rect 512958 433686 513014 433714
rect 513048 433714 513056 433720
rect 513090 433720 513156 433748
rect 513090 433714 513104 433720
rect 513048 433686 513104 433714
rect 513138 433714 513156 433720
rect 513190 433720 513256 433748
rect 513290 433720 513377 433748
rect 513190 433714 513194 433720
rect 513138 433686 513194 433714
rect 513228 433714 513256 433720
rect 513228 433686 513284 433714
rect 513318 433686 513377 433720
rect 512683 433627 513377 433686
rect 513439 434290 513458 434324
rect 513492 434308 513674 434324
rect 513492 434290 513605 434308
rect 513439 434274 513605 434290
rect 513639 434274 513674 434308
rect 513439 434234 513674 434274
rect 513439 434200 513458 434234
rect 513492 434218 513674 434234
rect 513492 434200 513605 434218
rect 513439 434184 513605 434200
rect 513639 434184 513674 434218
rect 513439 434144 513674 434184
rect 513439 434110 513458 434144
rect 513492 434128 513674 434144
rect 513492 434110 513605 434128
rect 513439 434094 513605 434110
rect 513639 434094 513674 434128
rect 513439 434054 513674 434094
rect 513439 434020 513458 434054
rect 513492 434038 513674 434054
rect 513492 434020 513605 434038
rect 513439 434004 513605 434020
rect 513639 434004 513674 434038
rect 513439 433964 513674 434004
rect 513439 433930 513458 433964
rect 513492 433948 513674 433964
rect 513492 433930 513605 433948
rect 513439 433914 513605 433930
rect 513639 433914 513674 433948
rect 513439 433874 513674 433914
rect 513439 433840 513458 433874
rect 513492 433858 513674 433874
rect 513492 433840 513605 433858
rect 513439 433824 513605 433840
rect 513639 433824 513674 433858
rect 513439 433784 513674 433824
rect 513439 433750 513458 433784
rect 513492 433768 513674 433784
rect 513492 433750 513605 433768
rect 513439 433734 513605 433750
rect 513639 433734 513674 433768
rect 513439 433694 513674 433734
rect 513439 433660 513458 433694
rect 513492 433678 513674 433694
rect 513492 433660 513605 433678
rect 513439 433644 513605 433660
rect 513639 433644 513674 433678
rect 512151 433570 512170 433604
rect 512204 433588 512621 433604
rect 512204 433570 512317 433588
rect 512151 433565 512317 433570
rect 511164 433554 512317 433565
rect 512351 433554 512418 433588
rect 512452 433565 512621 433588
rect 513439 433604 513674 433644
rect 513439 433570 513458 433604
rect 513492 433588 513674 433604
rect 513492 433570 513605 433588
rect 513439 433565 513605 433570
rect 512452 433554 513605 433565
rect 513639 433554 513674 433588
rect 503370 433546 513674 433554
rect 503370 433512 503646 433546
rect 503680 433512 503736 433546
rect 503770 433512 503826 433546
rect 503860 433512 503916 433546
rect 503950 433512 504006 433546
rect 504040 433512 504096 433546
rect 504130 433512 504186 433546
rect 504220 433512 504276 433546
rect 504310 433512 504366 433546
rect 504400 433512 504934 433546
rect 504968 433512 505024 433546
rect 505058 433512 505114 433546
rect 505148 433512 505204 433546
rect 505238 433512 505294 433546
rect 505328 433512 505384 433546
rect 505418 433512 505474 433546
rect 505508 433512 505564 433546
rect 505598 433512 505654 433546
rect 505688 433512 506222 433546
rect 506256 433512 506312 433546
rect 506346 433512 506402 433546
rect 506436 433512 506492 433546
rect 506526 433512 506582 433546
rect 506616 433512 506672 433546
rect 506706 433512 506762 433546
rect 506796 433512 506852 433546
rect 506886 433512 506942 433546
rect 506976 433512 507510 433546
rect 507544 433512 507600 433546
rect 507634 433512 507690 433546
rect 507724 433512 507780 433546
rect 507814 433512 507870 433546
rect 507904 433512 507960 433546
rect 507994 433512 508050 433546
rect 508084 433512 508140 433546
rect 508174 433512 508230 433546
rect 508264 433512 508798 433546
rect 508832 433512 508888 433546
rect 508922 433512 508978 433546
rect 509012 433512 509068 433546
rect 509102 433512 509158 433546
rect 509192 433512 509248 433546
rect 509282 433512 509338 433546
rect 509372 433512 509428 433546
rect 509462 433512 509518 433546
rect 509552 433512 510086 433546
rect 510120 433512 510176 433546
rect 510210 433512 510266 433546
rect 510300 433512 510356 433546
rect 510390 433512 510446 433546
rect 510480 433512 510536 433546
rect 510570 433512 510626 433546
rect 510660 433512 510716 433546
rect 510750 433512 510806 433546
rect 510840 433512 511374 433546
rect 511408 433512 511464 433546
rect 511498 433512 511554 433546
rect 511588 433512 511644 433546
rect 511678 433512 511734 433546
rect 511768 433512 511824 433546
rect 511858 433512 511914 433546
rect 511948 433512 512004 433546
rect 512038 433512 512094 433546
rect 512128 433512 512662 433546
rect 512696 433512 512752 433546
rect 512786 433512 512842 433546
rect 512876 433512 512932 433546
rect 512966 433512 513022 433546
rect 513056 433512 513112 433546
rect 513146 433512 513202 433546
rect 513236 433512 513292 433546
rect 513326 433512 513382 433546
rect 513416 433512 513674 433546
rect 503370 433498 513674 433512
rect 503370 433464 503402 433498
rect 503436 433464 504589 433498
rect 504623 433464 504690 433498
rect 504724 433464 505877 433498
rect 505911 433464 505978 433498
rect 506012 433464 507165 433498
rect 507199 433464 507266 433498
rect 507300 433464 508453 433498
rect 508487 433464 508554 433498
rect 508588 433464 509741 433498
rect 509775 433464 509842 433498
rect 509876 433464 511029 433498
rect 511063 433464 511130 433498
rect 511164 433464 512317 433498
rect 512351 433464 512418 433498
rect 512452 433464 513605 433498
rect 513639 433464 513674 433498
rect 501368 433284 501384 433408
rect 503370 433397 513674 433464
rect 503370 433363 503486 433397
rect 503520 433363 503576 433397
rect 503610 433363 503666 433397
rect 503700 433363 503756 433397
rect 503790 433363 503846 433397
rect 503880 433363 503936 433397
rect 503970 433363 504026 433397
rect 504060 433363 504116 433397
rect 504150 433363 504206 433397
rect 504240 433363 504296 433397
rect 504330 433363 504386 433397
rect 504420 433363 504476 433397
rect 504510 433363 504566 433397
rect 504600 433363 504774 433397
rect 504808 433363 504864 433397
rect 504898 433363 504954 433397
rect 504988 433363 505044 433397
rect 505078 433363 505134 433397
rect 505168 433363 505224 433397
rect 505258 433363 505314 433397
rect 505348 433363 505404 433397
rect 505438 433363 505494 433397
rect 505528 433363 505584 433397
rect 505618 433363 505674 433397
rect 505708 433363 505764 433397
rect 505798 433363 505854 433397
rect 505888 433363 506062 433397
rect 506096 433363 506152 433397
rect 506186 433363 506242 433397
rect 506276 433363 506332 433397
rect 506366 433363 506422 433397
rect 506456 433363 506512 433397
rect 506546 433363 506602 433397
rect 506636 433363 506692 433397
rect 506726 433363 506782 433397
rect 506816 433363 506872 433397
rect 506906 433363 506962 433397
rect 506996 433363 507052 433397
rect 507086 433363 507142 433397
rect 507176 433363 507350 433397
rect 507384 433363 507440 433397
rect 507474 433363 507530 433397
rect 507564 433363 507620 433397
rect 507654 433363 507710 433397
rect 507744 433363 507800 433397
rect 507834 433363 507890 433397
rect 507924 433363 507980 433397
rect 508014 433363 508070 433397
rect 508104 433363 508160 433397
rect 508194 433363 508250 433397
rect 508284 433363 508340 433397
rect 508374 433363 508430 433397
rect 508464 433363 508638 433397
rect 508672 433363 508728 433397
rect 508762 433363 508818 433397
rect 508852 433363 508908 433397
rect 508942 433363 508998 433397
rect 509032 433363 509088 433397
rect 509122 433363 509178 433397
rect 509212 433363 509268 433397
rect 509302 433363 509358 433397
rect 509392 433363 509448 433397
rect 509482 433363 509538 433397
rect 509572 433363 509628 433397
rect 509662 433363 509718 433397
rect 509752 433363 509926 433397
rect 509960 433363 510016 433397
rect 510050 433363 510106 433397
rect 510140 433363 510196 433397
rect 510230 433363 510286 433397
rect 510320 433363 510376 433397
rect 510410 433363 510466 433397
rect 510500 433363 510556 433397
rect 510590 433363 510646 433397
rect 510680 433363 510736 433397
rect 510770 433363 510826 433397
rect 510860 433363 510916 433397
rect 510950 433363 511006 433397
rect 511040 433363 511214 433397
rect 511248 433363 511304 433397
rect 511338 433363 511394 433397
rect 511428 433363 511484 433397
rect 511518 433363 511574 433397
rect 511608 433363 511664 433397
rect 511698 433363 511754 433397
rect 511788 433363 511844 433397
rect 511878 433363 511934 433397
rect 511968 433363 512024 433397
rect 512058 433363 512114 433397
rect 512148 433363 512204 433397
rect 512238 433363 512294 433397
rect 512328 433363 512502 433397
rect 512536 433363 512592 433397
rect 512626 433363 512682 433397
rect 512716 433363 512772 433397
rect 512806 433363 512862 433397
rect 512896 433363 512952 433397
rect 512986 433363 513042 433397
rect 513076 433363 513132 433397
rect 513166 433363 513222 433397
rect 513256 433363 513312 433397
rect 513346 433363 513402 433397
rect 513436 433363 513492 433397
rect 513526 433363 513582 433397
rect 513616 433363 513674 433397
rect 503370 433296 513674 433363
rect 503370 433262 503486 433296
rect 503520 433262 503576 433296
rect 503610 433262 503666 433296
rect 503700 433262 503756 433296
rect 503790 433262 503846 433296
rect 503880 433262 503936 433296
rect 503970 433262 504026 433296
rect 504060 433262 504116 433296
rect 504150 433262 504206 433296
rect 504240 433262 504296 433296
rect 504330 433262 504386 433296
rect 504420 433262 504476 433296
rect 504510 433262 504566 433296
rect 504600 433262 504774 433296
rect 504808 433262 504864 433296
rect 504898 433262 504954 433296
rect 504988 433262 505044 433296
rect 505078 433262 505134 433296
rect 505168 433262 505224 433296
rect 505258 433262 505314 433296
rect 505348 433262 505404 433296
rect 505438 433262 505494 433296
rect 505528 433262 505584 433296
rect 505618 433262 505674 433296
rect 505708 433262 505764 433296
rect 505798 433262 505854 433296
rect 505888 433262 506062 433296
rect 506096 433262 506152 433296
rect 506186 433262 506242 433296
rect 506276 433262 506332 433296
rect 506366 433262 506422 433296
rect 506456 433262 506512 433296
rect 506546 433262 506602 433296
rect 506636 433262 506692 433296
rect 506726 433262 506782 433296
rect 506816 433262 506872 433296
rect 506906 433262 506962 433296
rect 506996 433262 507052 433296
rect 507086 433262 507142 433296
rect 507176 433262 507350 433296
rect 507384 433262 507440 433296
rect 507474 433262 507530 433296
rect 507564 433262 507620 433296
rect 507654 433262 507710 433296
rect 507744 433262 507800 433296
rect 507834 433262 507890 433296
rect 507924 433262 507980 433296
rect 508014 433262 508070 433296
rect 508104 433262 508160 433296
rect 508194 433262 508250 433296
rect 508284 433262 508340 433296
rect 508374 433262 508430 433296
rect 508464 433262 508638 433296
rect 508672 433262 508728 433296
rect 508762 433262 508818 433296
rect 508852 433262 508908 433296
rect 508942 433262 508998 433296
rect 509032 433262 509088 433296
rect 509122 433262 509178 433296
rect 509212 433262 509268 433296
rect 509302 433262 509358 433296
rect 509392 433262 509448 433296
rect 509482 433262 509538 433296
rect 509572 433262 509628 433296
rect 509662 433262 509718 433296
rect 509752 433262 509926 433296
rect 509960 433262 510016 433296
rect 510050 433262 510106 433296
rect 510140 433262 510196 433296
rect 510230 433262 510286 433296
rect 510320 433262 510376 433296
rect 510410 433262 510466 433296
rect 510500 433262 510556 433296
rect 510590 433262 510646 433296
rect 510680 433262 510736 433296
rect 510770 433262 510826 433296
rect 510860 433262 510916 433296
rect 510950 433262 511006 433296
rect 511040 433262 511214 433296
rect 511248 433262 511304 433296
rect 511338 433262 511394 433296
rect 511428 433262 511484 433296
rect 511518 433262 511574 433296
rect 511608 433262 511664 433296
rect 511698 433262 511754 433296
rect 511788 433262 511844 433296
rect 511878 433262 511934 433296
rect 511968 433262 512024 433296
rect 512058 433262 512114 433296
rect 512148 433262 512204 433296
rect 512238 433262 512294 433296
rect 512328 433262 512502 433296
rect 512536 433262 512592 433296
rect 512626 433262 512682 433296
rect 512716 433262 512772 433296
rect 512806 433262 512862 433296
rect 512896 433262 512952 433296
rect 512986 433262 513042 433296
rect 513076 433262 513132 433296
rect 513166 433262 513222 433296
rect 513256 433262 513312 433296
rect 513346 433262 513402 433296
rect 513436 433262 513492 433296
rect 513526 433262 513582 433296
rect 513616 433262 513674 433296
rect 503370 433200 513674 433262
rect 501368 433060 501384 433184
rect 503370 433166 503402 433200
rect 503436 433166 504589 433200
rect 504623 433166 504690 433200
rect 504724 433166 505877 433200
rect 505911 433166 505978 433200
rect 506012 433166 507165 433200
rect 507199 433166 507266 433200
rect 507300 433166 508453 433200
rect 508487 433166 508554 433200
rect 508588 433166 509741 433200
rect 509775 433166 509842 433200
rect 509876 433166 511029 433200
rect 511063 433166 511130 433200
rect 511164 433166 512317 433200
rect 512351 433166 512418 433200
rect 512452 433166 513605 433200
rect 513639 433166 513674 433200
rect 503370 433148 513674 433166
rect 503370 433114 503665 433148
rect 503699 433114 503755 433148
rect 503789 433114 503845 433148
rect 503879 433114 503935 433148
rect 503969 433114 504025 433148
rect 504059 433114 504115 433148
rect 504149 433114 504205 433148
rect 504239 433114 504295 433148
rect 504329 433114 504385 433148
rect 504419 433114 504953 433148
rect 504987 433114 505043 433148
rect 505077 433114 505133 433148
rect 505167 433114 505223 433148
rect 505257 433114 505313 433148
rect 505347 433114 505403 433148
rect 505437 433114 505493 433148
rect 505527 433114 505583 433148
rect 505617 433114 505673 433148
rect 505707 433114 506241 433148
rect 506275 433114 506331 433148
rect 506365 433114 506421 433148
rect 506455 433114 506511 433148
rect 506545 433114 506601 433148
rect 506635 433114 506691 433148
rect 506725 433114 506781 433148
rect 506815 433114 506871 433148
rect 506905 433114 506961 433148
rect 506995 433114 507529 433148
rect 507563 433114 507619 433148
rect 507653 433114 507709 433148
rect 507743 433114 507799 433148
rect 507833 433114 507889 433148
rect 507923 433114 507979 433148
rect 508013 433114 508069 433148
rect 508103 433114 508159 433148
rect 508193 433114 508249 433148
rect 508283 433114 508817 433148
rect 508851 433114 508907 433148
rect 508941 433114 508997 433148
rect 509031 433114 509087 433148
rect 509121 433114 509177 433148
rect 509211 433114 509267 433148
rect 509301 433114 509357 433148
rect 509391 433114 509447 433148
rect 509481 433114 509537 433148
rect 509571 433114 510105 433148
rect 510139 433114 510195 433148
rect 510229 433114 510285 433148
rect 510319 433114 510375 433148
rect 510409 433114 510465 433148
rect 510499 433114 510555 433148
rect 510589 433114 510645 433148
rect 510679 433114 510735 433148
rect 510769 433114 510825 433148
rect 510859 433114 511393 433148
rect 511427 433114 511483 433148
rect 511517 433114 511573 433148
rect 511607 433114 511663 433148
rect 511697 433114 511753 433148
rect 511787 433114 511843 433148
rect 511877 433114 511933 433148
rect 511967 433114 512023 433148
rect 512057 433114 512113 433148
rect 512147 433114 512681 433148
rect 512715 433114 512771 433148
rect 512805 433114 512861 433148
rect 512895 433114 512951 433148
rect 512985 433114 513041 433148
rect 513075 433114 513131 433148
rect 513165 433114 513221 433148
rect 513255 433114 513311 433148
rect 513345 433114 513401 433148
rect 513435 433114 513674 433148
rect 503370 433110 513674 433114
rect 503370 433076 503402 433110
rect 503436 433095 504589 433110
rect 503436 433076 503605 433095
rect 503370 433070 503605 433076
rect 500320 432068 500368 433044
rect 503370 433036 503552 433070
rect 503586 433036 503605 433070
rect 503370 433020 503605 433036
rect 504423 433076 504589 433095
rect 504623 433076 504690 433110
rect 504724 433095 505877 433110
rect 504724 433076 504893 433095
rect 504423 433070 504893 433076
rect 504423 433036 504840 433070
rect 504874 433036 504893 433070
rect 503370 432986 503402 433020
rect 503436 432986 503605 433020
rect 503370 432980 503605 432986
rect 501368 432836 501384 432960
rect 503370 432946 503552 432980
rect 503586 432946 503605 432980
rect 503370 432930 503605 432946
rect 503370 432896 503402 432930
rect 503436 432896 503605 432930
rect 503370 432890 503605 432896
rect 503370 432856 503552 432890
rect 503586 432856 503605 432890
rect 503370 432840 503605 432856
rect 503370 432806 503402 432840
rect 503436 432806 503605 432840
rect 503370 432800 503605 432806
rect 503370 432766 503552 432800
rect 503586 432766 503605 432800
rect 503370 432750 503605 432766
rect 501368 432612 501384 432736
rect 503370 432716 503402 432750
rect 503436 432716 503605 432750
rect 503370 432710 503605 432716
rect 503370 432676 503552 432710
rect 503586 432676 503605 432710
rect 503370 432660 503605 432676
rect 503370 432626 503402 432660
rect 503436 432626 503605 432660
rect 503370 432620 503605 432626
rect 503370 432586 503552 432620
rect 503586 432586 503605 432620
rect 503370 432570 503605 432586
rect 503370 432536 503402 432570
rect 503436 432536 503605 432570
rect 503370 432530 503605 432536
rect 501368 432388 501384 432512
rect 503370 432496 503552 432530
rect 503586 432496 503605 432530
rect 503370 432480 503605 432496
rect 503370 432446 503402 432480
rect 503436 432446 503605 432480
rect 503370 432440 503605 432446
rect 503370 432406 503552 432440
rect 503586 432406 503605 432440
rect 503370 432390 503605 432406
rect 503370 432356 503402 432390
rect 503436 432356 503605 432390
rect 503370 432350 503605 432356
rect 503370 432316 503552 432350
rect 503586 432316 503605 432350
rect 503667 432972 504361 433033
rect 503667 432938 503728 432972
rect 503762 432960 503818 432972
rect 503852 432960 503908 432972
rect 503942 432960 503998 432972
rect 503774 432938 503818 432960
rect 503874 432938 503908 432960
rect 503974 432938 503998 432960
rect 504032 432960 504088 432972
rect 504032 432938 504040 432960
rect 503667 432926 503740 432938
rect 503774 432926 503840 432938
rect 503874 432926 503940 432938
rect 503974 432926 504040 432938
rect 504074 432938 504088 432960
rect 504122 432960 504178 432972
rect 504122 432938 504140 432960
rect 504074 432926 504140 432938
rect 504174 432938 504178 432960
rect 504212 432960 504268 432972
rect 504212 432938 504240 432960
rect 504302 432938 504361 432972
rect 504174 432926 504240 432938
rect 504274 432926 504361 432938
rect 503667 432882 504361 432926
rect 503667 432848 503728 432882
rect 503762 432860 503818 432882
rect 503852 432860 503908 432882
rect 503942 432860 503998 432882
rect 503774 432848 503818 432860
rect 503874 432848 503908 432860
rect 503974 432848 503998 432860
rect 504032 432860 504088 432882
rect 504032 432848 504040 432860
rect 503667 432826 503740 432848
rect 503774 432826 503840 432848
rect 503874 432826 503940 432848
rect 503974 432826 504040 432848
rect 504074 432848 504088 432860
rect 504122 432860 504178 432882
rect 504122 432848 504140 432860
rect 504074 432826 504140 432848
rect 504174 432848 504178 432860
rect 504212 432860 504268 432882
rect 504212 432848 504240 432860
rect 504302 432848 504361 432882
rect 504174 432826 504240 432848
rect 504274 432826 504361 432848
rect 503667 432792 504361 432826
rect 503667 432758 503728 432792
rect 503762 432760 503818 432792
rect 503852 432760 503908 432792
rect 503942 432760 503998 432792
rect 503774 432758 503818 432760
rect 503874 432758 503908 432760
rect 503974 432758 503998 432760
rect 504032 432760 504088 432792
rect 504032 432758 504040 432760
rect 503667 432726 503740 432758
rect 503774 432726 503840 432758
rect 503874 432726 503940 432758
rect 503974 432726 504040 432758
rect 504074 432758 504088 432760
rect 504122 432760 504178 432792
rect 504122 432758 504140 432760
rect 504074 432726 504140 432758
rect 504174 432758 504178 432760
rect 504212 432760 504268 432792
rect 504212 432758 504240 432760
rect 504302 432758 504361 432792
rect 504174 432726 504240 432758
rect 504274 432726 504361 432758
rect 503667 432702 504361 432726
rect 503667 432668 503728 432702
rect 503762 432668 503818 432702
rect 503852 432668 503908 432702
rect 503942 432668 503998 432702
rect 504032 432668 504088 432702
rect 504122 432668 504178 432702
rect 504212 432668 504268 432702
rect 504302 432668 504361 432702
rect 503667 432660 504361 432668
rect 503667 432626 503740 432660
rect 503774 432626 503840 432660
rect 503874 432626 503940 432660
rect 503974 432626 504040 432660
rect 504074 432626 504140 432660
rect 504174 432626 504240 432660
rect 504274 432626 504361 432660
rect 503667 432612 504361 432626
rect 503667 432578 503728 432612
rect 503762 432578 503818 432612
rect 503852 432578 503908 432612
rect 503942 432578 503998 432612
rect 504032 432578 504088 432612
rect 504122 432578 504178 432612
rect 504212 432578 504268 432612
rect 504302 432578 504361 432612
rect 503667 432560 504361 432578
rect 503667 432526 503740 432560
rect 503774 432526 503840 432560
rect 503874 432526 503940 432560
rect 503974 432526 504040 432560
rect 504074 432526 504140 432560
rect 504174 432526 504240 432560
rect 504274 432526 504361 432560
rect 503667 432522 504361 432526
rect 503667 432488 503728 432522
rect 503762 432488 503818 432522
rect 503852 432488 503908 432522
rect 503942 432488 503998 432522
rect 504032 432488 504088 432522
rect 504122 432488 504178 432522
rect 504212 432488 504268 432522
rect 504302 432488 504361 432522
rect 503667 432460 504361 432488
rect 503667 432432 503740 432460
rect 503774 432432 503840 432460
rect 503874 432432 503940 432460
rect 503974 432432 504040 432460
rect 503667 432398 503728 432432
rect 503774 432426 503818 432432
rect 503874 432426 503908 432432
rect 503974 432426 503998 432432
rect 503762 432398 503818 432426
rect 503852 432398 503908 432426
rect 503942 432398 503998 432426
rect 504032 432426 504040 432432
rect 504074 432432 504140 432460
rect 504074 432426 504088 432432
rect 504032 432398 504088 432426
rect 504122 432426 504140 432432
rect 504174 432432 504240 432460
rect 504274 432432 504361 432460
rect 504174 432426 504178 432432
rect 504122 432398 504178 432426
rect 504212 432426 504240 432432
rect 504212 432398 504268 432426
rect 504302 432398 504361 432432
rect 503667 432339 504361 432398
rect 504423 433002 504442 433036
rect 504476 433020 504893 433036
rect 505711 433076 505877 433095
rect 505911 433076 505978 433110
rect 506012 433095 507165 433110
rect 506012 433076 506181 433095
rect 505711 433070 506181 433076
rect 505711 433036 506128 433070
rect 506162 433036 506181 433070
rect 504476 433002 504589 433020
rect 504423 432986 504589 433002
rect 504623 432986 504690 433020
rect 504724 432986 504893 433020
rect 504423 432980 504893 432986
rect 504423 432946 504840 432980
rect 504874 432946 504893 432980
rect 504423 432912 504442 432946
rect 504476 432930 504893 432946
rect 504476 432912 504589 432930
rect 504423 432896 504589 432912
rect 504623 432896 504690 432930
rect 504724 432896 504893 432930
rect 504423 432890 504893 432896
rect 504423 432856 504840 432890
rect 504874 432856 504893 432890
rect 504423 432822 504442 432856
rect 504476 432840 504893 432856
rect 504476 432822 504589 432840
rect 504423 432806 504589 432822
rect 504623 432806 504690 432840
rect 504724 432806 504893 432840
rect 504423 432800 504893 432806
rect 504423 432766 504840 432800
rect 504874 432766 504893 432800
rect 504423 432732 504442 432766
rect 504476 432750 504893 432766
rect 504476 432732 504589 432750
rect 504423 432716 504589 432732
rect 504623 432716 504690 432750
rect 504724 432716 504893 432750
rect 504423 432710 504893 432716
rect 504423 432676 504840 432710
rect 504874 432676 504893 432710
rect 504423 432642 504442 432676
rect 504476 432660 504893 432676
rect 504476 432642 504589 432660
rect 504423 432626 504589 432642
rect 504623 432626 504690 432660
rect 504724 432626 504893 432660
rect 504423 432620 504893 432626
rect 504423 432586 504840 432620
rect 504874 432586 504893 432620
rect 504423 432552 504442 432586
rect 504476 432570 504893 432586
rect 504476 432552 504589 432570
rect 504423 432536 504589 432552
rect 504623 432536 504690 432570
rect 504724 432536 504893 432570
rect 504423 432530 504893 432536
rect 504423 432496 504840 432530
rect 504874 432496 504893 432530
rect 504423 432462 504442 432496
rect 504476 432480 504893 432496
rect 504476 432462 504589 432480
rect 504423 432446 504589 432462
rect 504623 432446 504690 432480
rect 504724 432446 504893 432480
rect 504423 432440 504893 432446
rect 504423 432406 504840 432440
rect 504874 432406 504893 432440
rect 504423 432372 504442 432406
rect 504476 432390 504893 432406
rect 504476 432372 504589 432390
rect 504423 432356 504589 432372
rect 504623 432356 504690 432390
rect 504724 432356 504893 432390
rect 504423 432350 504893 432356
rect 503370 432300 503605 432316
rect 501368 432164 501384 432288
rect 503370 432266 503402 432300
rect 503436 432277 503605 432300
rect 504423 432316 504840 432350
rect 504874 432316 504893 432350
rect 504955 432972 505649 433033
rect 504955 432938 505016 432972
rect 505050 432960 505106 432972
rect 505140 432960 505196 432972
rect 505230 432960 505286 432972
rect 505062 432938 505106 432960
rect 505162 432938 505196 432960
rect 505262 432938 505286 432960
rect 505320 432960 505376 432972
rect 505320 432938 505328 432960
rect 504955 432926 505028 432938
rect 505062 432926 505128 432938
rect 505162 432926 505228 432938
rect 505262 432926 505328 432938
rect 505362 432938 505376 432960
rect 505410 432960 505466 432972
rect 505410 432938 505428 432960
rect 505362 432926 505428 432938
rect 505462 432938 505466 432960
rect 505500 432960 505556 432972
rect 505500 432938 505528 432960
rect 505590 432938 505649 432972
rect 505462 432926 505528 432938
rect 505562 432926 505649 432938
rect 504955 432882 505649 432926
rect 504955 432848 505016 432882
rect 505050 432860 505106 432882
rect 505140 432860 505196 432882
rect 505230 432860 505286 432882
rect 505062 432848 505106 432860
rect 505162 432848 505196 432860
rect 505262 432848 505286 432860
rect 505320 432860 505376 432882
rect 505320 432848 505328 432860
rect 504955 432826 505028 432848
rect 505062 432826 505128 432848
rect 505162 432826 505228 432848
rect 505262 432826 505328 432848
rect 505362 432848 505376 432860
rect 505410 432860 505466 432882
rect 505410 432848 505428 432860
rect 505362 432826 505428 432848
rect 505462 432848 505466 432860
rect 505500 432860 505556 432882
rect 505500 432848 505528 432860
rect 505590 432848 505649 432882
rect 505462 432826 505528 432848
rect 505562 432826 505649 432848
rect 504955 432792 505649 432826
rect 504955 432758 505016 432792
rect 505050 432760 505106 432792
rect 505140 432760 505196 432792
rect 505230 432760 505286 432792
rect 505062 432758 505106 432760
rect 505162 432758 505196 432760
rect 505262 432758 505286 432760
rect 505320 432760 505376 432792
rect 505320 432758 505328 432760
rect 504955 432726 505028 432758
rect 505062 432726 505128 432758
rect 505162 432726 505228 432758
rect 505262 432726 505328 432758
rect 505362 432758 505376 432760
rect 505410 432760 505466 432792
rect 505410 432758 505428 432760
rect 505362 432726 505428 432758
rect 505462 432758 505466 432760
rect 505500 432760 505556 432792
rect 505500 432758 505528 432760
rect 505590 432758 505649 432792
rect 505462 432726 505528 432758
rect 505562 432726 505649 432758
rect 504955 432702 505649 432726
rect 504955 432668 505016 432702
rect 505050 432668 505106 432702
rect 505140 432668 505196 432702
rect 505230 432668 505286 432702
rect 505320 432668 505376 432702
rect 505410 432668 505466 432702
rect 505500 432668 505556 432702
rect 505590 432668 505649 432702
rect 504955 432660 505649 432668
rect 504955 432626 505028 432660
rect 505062 432626 505128 432660
rect 505162 432626 505228 432660
rect 505262 432626 505328 432660
rect 505362 432626 505428 432660
rect 505462 432626 505528 432660
rect 505562 432626 505649 432660
rect 504955 432612 505649 432626
rect 504955 432578 505016 432612
rect 505050 432578 505106 432612
rect 505140 432578 505196 432612
rect 505230 432578 505286 432612
rect 505320 432578 505376 432612
rect 505410 432578 505466 432612
rect 505500 432578 505556 432612
rect 505590 432578 505649 432612
rect 504955 432560 505649 432578
rect 504955 432526 505028 432560
rect 505062 432526 505128 432560
rect 505162 432526 505228 432560
rect 505262 432526 505328 432560
rect 505362 432526 505428 432560
rect 505462 432526 505528 432560
rect 505562 432526 505649 432560
rect 504955 432522 505649 432526
rect 504955 432488 505016 432522
rect 505050 432488 505106 432522
rect 505140 432488 505196 432522
rect 505230 432488 505286 432522
rect 505320 432488 505376 432522
rect 505410 432488 505466 432522
rect 505500 432488 505556 432522
rect 505590 432488 505649 432522
rect 504955 432460 505649 432488
rect 504955 432432 505028 432460
rect 505062 432432 505128 432460
rect 505162 432432 505228 432460
rect 505262 432432 505328 432460
rect 504955 432398 505016 432432
rect 505062 432426 505106 432432
rect 505162 432426 505196 432432
rect 505262 432426 505286 432432
rect 505050 432398 505106 432426
rect 505140 432398 505196 432426
rect 505230 432398 505286 432426
rect 505320 432426 505328 432432
rect 505362 432432 505428 432460
rect 505362 432426 505376 432432
rect 505320 432398 505376 432426
rect 505410 432426 505428 432432
rect 505462 432432 505528 432460
rect 505562 432432 505649 432460
rect 505462 432426 505466 432432
rect 505410 432398 505466 432426
rect 505500 432426 505528 432432
rect 505500 432398 505556 432426
rect 505590 432398 505649 432432
rect 504955 432339 505649 432398
rect 505711 433002 505730 433036
rect 505764 433020 506181 433036
rect 506999 433076 507165 433095
rect 507199 433076 507266 433110
rect 507300 433095 508453 433110
rect 507300 433076 507469 433095
rect 506999 433070 507469 433076
rect 506999 433036 507416 433070
rect 507450 433036 507469 433070
rect 505764 433002 505877 433020
rect 505711 432986 505877 433002
rect 505911 432986 505978 433020
rect 506012 432986 506181 433020
rect 505711 432980 506181 432986
rect 505711 432946 506128 432980
rect 506162 432946 506181 432980
rect 505711 432912 505730 432946
rect 505764 432930 506181 432946
rect 505764 432912 505877 432930
rect 505711 432896 505877 432912
rect 505911 432896 505978 432930
rect 506012 432896 506181 432930
rect 505711 432890 506181 432896
rect 505711 432856 506128 432890
rect 506162 432856 506181 432890
rect 505711 432822 505730 432856
rect 505764 432840 506181 432856
rect 505764 432822 505877 432840
rect 505711 432806 505877 432822
rect 505911 432806 505978 432840
rect 506012 432806 506181 432840
rect 505711 432800 506181 432806
rect 505711 432766 506128 432800
rect 506162 432766 506181 432800
rect 505711 432732 505730 432766
rect 505764 432750 506181 432766
rect 505764 432732 505877 432750
rect 505711 432716 505877 432732
rect 505911 432716 505978 432750
rect 506012 432716 506181 432750
rect 505711 432710 506181 432716
rect 505711 432676 506128 432710
rect 506162 432676 506181 432710
rect 505711 432642 505730 432676
rect 505764 432660 506181 432676
rect 505764 432642 505877 432660
rect 505711 432626 505877 432642
rect 505911 432626 505978 432660
rect 506012 432626 506181 432660
rect 505711 432620 506181 432626
rect 505711 432586 506128 432620
rect 506162 432586 506181 432620
rect 505711 432552 505730 432586
rect 505764 432570 506181 432586
rect 505764 432552 505877 432570
rect 505711 432536 505877 432552
rect 505911 432536 505978 432570
rect 506012 432536 506181 432570
rect 505711 432530 506181 432536
rect 505711 432496 506128 432530
rect 506162 432496 506181 432530
rect 505711 432462 505730 432496
rect 505764 432480 506181 432496
rect 505764 432462 505877 432480
rect 505711 432446 505877 432462
rect 505911 432446 505978 432480
rect 506012 432446 506181 432480
rect 505711 432440 506181 432446
rect 505711 432406 506128 432440
rect 506162 432406 506181 432440
rect 505711 432372 505730 432406
rect 505764 432390 506181 432406
rect 505764 432372 505877 432390
rect 505711 432356 505877 432372
rect 505911 432356 505978 432390
rect 506012 432356 506181 432390
rect 505711 432350 506181 432356
rect 504423 432282 504442 432316
rect 504476 432300 504893 432316
rect 504476 432282 504589 432300
rect 504423 432277 504589 432282
rect 503436 432266 504589 432277
rect 504623 432266 504690 432300
rect 504724 432277 504893 432300
rect 505711 432316 506128 432350
rect 506162 432316 506181 432350
rect 506243 432972 506937 433033
rect 506243 432938 506304 432972
rect 506338 432960 506394 432972
rect 506428 432960 506484 432972
rect 506518 432960 506574 432972
rect 506350 432938 506394 432960
rect 506450 432938 506484 432960
rect 506550 432938 506574 432960
rect 506608 432960 506664 432972
rect 506608 432938 506616 432960
rect 506243 432926 506316 432938
rect 506350 432926 506416 432938
rect 506450 432926 506516 432938
rect 506550 432926 506616 432938
rect 506650 432938 506664 432960
rect 506698 432960 506754 432972
rect 506698 432938 506716 432960
rect 506650 432926 506716 432938
rect 506750 432938 506754 432960
rect 506788 432960 506844 432972
rect 506788 432938 506816 432960
rect 506878 432938 506937 432972
rect 506750 432926 506816 432938
rect 506850 432926 506937 432938
rect 506243 432882 506937 432926
rect 506243 432848 506304 432882
rect 506338 432860 506394 432882
rect 506428 432860 506484 432882
rect 506518 432860 506574 432882
rect 506350 432848 506394 432860
rect 506450 432848 506484 432860
rect 506550 432848 506574 432860
rect 506608 432860 506664 432882
rect 506608 432848 506616 432860
rect 506243 432826 506316 432848
rect 506350 432826 506416 432848
rect 506450 432826 506516 432848
rect 506550 432826 506616 432848
rect 506650 432848 506664 432860
rect 506698 432860 506754 432882
rect 506698 432848 506716 432860
rect 506650 432826 506716 432848
rect 506750 432848 506754 432860
rect 506788 432860 506844 432882
rect 506788 432848 506816 432860
rect 506878 432848 506937 432882
rect 506750 432826 506816 432848
rect 506850 432826 506937 432848
rect 506243 432792 506937 432826
rect 506243 432758 506304 432792
rect 506338 432760 506394 432792
rect 506428 432760 506484 432792
rect 506518 432760 506574 432792
rect 506350 432758 506394 432760
rect 506450 432758 506484 432760
rect 506550 432758 506574 432760
rect 506608 432760 506664 432792
rect 506608 432758 506616 432760
rect 506243 432726 506316 432758
rect 506350 432726 506416 432758
rect 506450 432726 506516 432758
rect 506550 432726 506616 432758
rect 506650 432758 506664 432760
rect 506698 432760 506754 432792
rect 506698 432758 506716 432760
rect 506650 432726 506716 432758
rect 506750 432758 506754 432760
rect 506788 432760 506844 432792
rect 506788 432758 506816 432760
rect 506878 432758 506937 432792
rect 506750 432726 506816 432758
rect 506850 432726 506937 432758
rect 506243 432702 506937 432726
rect 506243 432668 506304 432702
rect 506338 432668 506394 432702
rect 506428 432668 506484 432702
rect 506518 432668 506574 432702
rect 506608 432668 506664 432702
rect 506698 432668 506754 432702
rect 506788 432668 506844 432702
rect 506878 432668 506937 432702
rect 506243 432660 506937 432668
rect 506243 432626 506316 432660
rect 506350 432626 506416 432660
rect 506450 432626 506516 432660
rect 506550 432626 506616 432660
rect 506650 432626 506716 432660
rect 506750 432626 506816 432660
rect 506850 432626 506937 432660
rect 506243 432612 506937 432626
rect 506243 432578 506304 432612
rect 506338 432578 506394 432612
rect 506428 432578 506484 432612
rect 506518 432578 506574 432612
rect 506608 432578 506664 432612
rect 506698 432578 506754 432612
rect 506788 432578 506844 432612
rect 506878 432578 506937 432612
rect 506243 432560 506937 432578
rect 506243 432526 506316 432560
rect 506350 432526 506416 432560
rect 506450 432526 506516 432560
rect 506550 432526 506616 432560
rect 506650 432526 506716 432560
rect 506750 432526 506816 432560
rect 506850 432526 506937 432560
rect 506243 432522 506937 432526
rect 506243 432488 506304 432522
rect 506338 432488 506394 432522
rect 506428 432488 506484 432522
rect 506518 432488 506574 432522
rect 506608 432488 506664 432522
rect 506698 432488 506754 432522
rect 506788 432488 506844 432522
rect 506878 432488 506937 432522
rect 506243 432460 506937 432488
rect 506243 432432 506316 432460
rect 506350 432432 506416 432460
rect 506450 432432 506516 432460
rect 506550 432432 506616 432460
rect 506243 432398 506304 432432
rect 506350 432426 506394 432432
rect 506450 432426 506484 432432
rect 506550 432426 506574 432432
rect 506338 432398 506394 432426
rect 506428 432398 506484 432426
rect 506518 432398 506574 432426
rect 506608 432426 506616 432432
rect 506650 432432 506716 432460
rect 506650 432426 506664 432432
rect 506608 432398 506664 432426
rect 506698 432426 506716 432432
rect 506750 432432 506816 432460
rect 506850 432432 506937 432460
rect 506750 432426 506754 432432
rect 506698 432398 506754 432426
rect 506788 432426 506816 432432
rect 506788 432398 506844 432426
rect 506878 432398 506937 432432
rect 506243 432339 506937 432398
rect 506999 433002 507018 433036
rect 507052 433020 507469 433036
rect 508287 433076 508453 433095
rect 508487 433076 508554 433110
rect 508588 433095 509741 433110
rect 508588 433076 508757 433095
rect 508287 433070 508757 433076
rect 508287 433036 508704 433070
rect 508738 433036 508757 433070
rect 507052 433002 507165 433020
rect 506999 432986 507165 433002
rect 507199 432986 507266 433020
rect 507300 432986 507469 433020
rect 506999 432980 507469 432986
rect 506999 432946 507416 432980
rect 507450 432946 507469 432980
rect 506999 432912 507018 432946
rect 507052 432930 507469 432946
rect 507052 432912 507165 432930
rect 506999 432896 507165 432912
rect 507199 432896 507266 432930
rect 507300 432896 507469 432930
rect 506999 432890 507469 432896
rect 506999 432856 507416 432890
rect 507450 432856 507469 432890
rect 506999 432822 507018 432856
rect 507052 432840 507469 432856
rect 507052 432822 507165 432840
rect 506999 432806 507165 432822
rect 507199 432806 507266 432840
rect 507300 432806 507469 432840
rect 506999 432800 507469 432806
rect 506999 432766 507416 432800
rect 507450 432766 507469 432800
rect 506999 432732 507018 432766
rect 507052 432750 507469 432766
rect 507052 432732 507165 432750
rect 506999 432716 507165 432732
rect 507199 432716 507266 432750
rect 507300 432716 507469 432750
rect 506999 432710 507469 432716
rect 506999 432676 507416 432710
rect 507450 432676 507469 432710
rect 506999 432642 507018 432676
rect 507052 432660 507469 432676
rect 507052 432642 507165 432660
rect 506999 432626 507165 432642
rect 507199 432626 507266 432660
rect 507300 432626 507469 432660
rect 506999 432620 507469 432626
rect 506999 432586 507416 432620
rect 507450 432586 507469 432620
rect 506999 432552 507018 432586
rect 507052 432570 507469 432586
rect 507052 432552 507165 432570
rect 506999 432536 507165 432552
rect 507199 432536 507266 432570
rect 507300 432536 507469 432570
rect 506999 432530 507469 432536
rect 506999 432496 507416 432530
rect 507450 432496 507469 432530
rect 506999 432462 507018 432496
rect 507052 432480 507469 432496
rect 507052 432462 507165 432480
rect 506999 432446 507165 432462
rect 507199 432446 507266 432480
rect 507300 432446 507469 432480
rect 506999 432440 507469 432446
rect 506999 432406 507416 432440
rect 507450 432406 507469 432440
rect 506999 432372 507018 432406
rect 507052 432390 507469 432406
rect 507052 432372 507165 432390
rect 506999 432356 507165 432372
rect 507199 432356 507266 432390
rect 507300 432356 507469 432390
rect 506999 432350 507469 432356
rect 505711 432282 505730 432316
rect 505764 432300 506181 432316
rect 505764 432282 505877 432300
rect 505711 432277 505877 432282
rect 504724 432266 505877 432277
rect 505911 432266 505978 432300
rect 506012 432277 506181 432300
rect 506999 432316 507416 432350
rect 507450 432316 507469 432350
rect 507531 432972 508225 433033
rect 507531 432938 507592 432972
rect 507626 432960 507682 432972
rect 507716 432960 507772 432972
rect 507806 432960 507862 432972
rect 507638 432938 507682 432960
rect 507738 432938 507772 432960
rect 507838 432938 507862 432960
rect 507896 432960 507952 432972
rect 507896 432938 507904 432960
rect 507531 432926 507604 432938
rect 507638 432926 507704 432938
rect 507738 432926 507804 432938
rect 507838 432926 507904 432938
rect 507938 432938 507952 432960
rect 507986 432960 508042 432972
rect 507986 432938 508004 432960
rect 507938 432926 508004 432938
rect 508038 432938 508042 432960
rect 508076 432960 508132 432972
rect 508076 432938 508104 432960
rect 508166 432938 508225 432972
rect 508038 432926 508104 432938
rect 508138 432926 508225 432938
rect 507531 432882 508225 432926
rect 507531 432848 507592 432882
rect 507626 432860 507682 432882
rect 507716 432860 507772 432882
rect 507806 432860 507862 432882
rect 507638 432848 507682 432860
rect 507738 432848 507772 432860
rect 507838 432848 507862 432860
rect 507896 432860 507952 432882
rect 507896 432848 507904 432860
rect 507531 432826 507604 432848
rect 507638 432826 507704 432848
rect 507738 432826 507804 432848
rect 507838 432826 507904 432848
rect 507938 432848 507952 432860
rect 507986 432860 508042 432882
rect 507986 432848 508004 432860
rect 507938 432826 508004 432848
rect 508038 432848 508042 432860
rect 508076 432860 508132 432882
rect 508076 432848 508104 432860
rect 508166 432848 508225 432882
rect 508038 432826 508104 432848
rect 508138 432826 508225 432848
rect 507531 432792 508225 432826
rect 507531 432758 507592 432792
rect 507626 432760 507682 432792
rect 507716 432760 507772 432792
rect 507806 432760 507862 432792
rect 507638 432758 507682 432760
rect 507738 432758 507772 432760
rect 507838 432758 507862 432760
rect 507896 432760 507952 432792
rect 507896 432758 507904 432760
rect 507531 432726 507604 432758
rect 507638 432726 507704 432758
rect 507738 432726 507804 432758
rect 507838 432726 507904 432758
rect 507938 432758 507952 432760
rect 507986 432760 508042 432792
rect 507986 432758 508004 432760
rect 507938 432726 508004 432758
rect 508038 432758 508042 432760
rect 508076 432760 508132 432792
rect 508076 432758 508104 432760
rect 508166 432758 508225 432792
rect 508038 432726 508104 432758
rect 508138 432726 508225 432758
rect 507531 432702 508225 432726
rect 507531 432668 507592 432702
rect 507626 432668 507682 432702
rect 507716 432668 507772 432702
rect 507806 432668 507862 432702
rect 507896 432668 507952 432702
rect 507986 432668 508042 432702
rect 508076 432668 508132 432702
rect 508166 432668 508225 432702
rect 507531 432660 508225 432668
rect 507531 432626 507604 432660
rect 507638 432626 507704 432660
rect 507738 432626 507804 432660
rect 507838 432626 507904 432660
rect 507938 432626 508004 432660
rect 508038 432626 508104 432660
rect 508138 432626 508225 432660
rect 507531 432612 508225 432626
rect 507531 432578 507592 432612
rect 507626 432578 507682 432612
rect 507716 432578 507772 432612
rect 507806 432578 507862 432612
rect 507896 432578 507952 432612
rect 507986 432578 508042 432612
rect 508076 432578 508132 432612
rect 508166 432578 508225 432612
rect 507531 432560 508225 432578
rect 507531 432526 507604 432560
rect 507638 432526 507704 432560
rect 507738 432526 507804 432560
rect 507838 432526 507904 432560
rect 507938 432526 508004 432560
rect 508038 432526 508104 432560
rect 508138 432526 508225 432560
rect 507531 432522 508225 432526
rect 507531 432488 507592 432522
rect 507626 432488 507682 432522
rect 507716 432488 507772 432522
rect 507806 432488 507862 432522
rect 507896 432488 507952 432522
rect 507986 432488 508042 432522
rect 508076 432488 508132 432522
rect 508166 432488 508225 432522
rect 507531 432460 508225 432488
rect 507531 432432 507604 432460
rect 507638 432432 507704 432460
rect 507738 432432 507804 432460
rect 507838 432432 507904 432460
rect 507531 432398 507592 432432
rect 507638 432426 507682 432432
rect 507738 432426 507772 432432
rect 507838 432426 507862 432432
rect 507626 432398 507682 432426
rect 507716 432398 507772 432426
rect 507806 432398 507862 432426
rect 507896 432426 507904 432432
rect 507938 432432 508004 432460
rect 507938 432426 507952 432432
rect 507896 432398 507952 432426
rect 507986 432426 508004 432432
rect 508038 432432 508104 432460
rect 508138 432432 508225 432460
rect 508038 432426 508042 432432
rect 507986 432398 508042 432426
rect 508076 432426 508104 432432
rect 508076 432398 508132 432426
rect 508166 432398 508225 432432
rect 507531 432339 508225 432398
rect 508287 433002 508306 433036
rect 508340 433020 508757 433036
rect 509575 433076 509741 433095
rect 509775 433076 509842 433110
rect 509876 433095 511029 433110
rect 509876 433076 510045 433095
rect 509575 433070 510045 433076
rect 509575 433036 509992 433070
rect 510026 433036 510045 433070
rect 508340 433002 508453 433020
rect 508287 432986 508453 433002
rect 508487 432986 508554 433020
rect 508588 432986 508757 433020
rect 508287 432980 508757 432986
rect 508287 432946 508704 432980
rect 508738 432946 508757 432980
rect 508287 432912 508306 432946
rect 508340 432930 508757 432946
rect 508340 432912 508453 432930
rect 508287 432896 508453 432912
rect 508487 432896 508554 432930
rect 508588 432896 508757 432930
rect 508287 432890 508757 432896
rect 508287 432856 508704 432890
rect 508738 432856 508757 432890
rect 508287 432822 508306 432856
rect 508340 432840 508757 432856
rect 508340 432822 508453 432840
rect 508287 432806 508453 432822
rect 508487 432806 508554 432840
rect 508588 432806 508757 432840
rect 508287 432800 508757 432806
rect 508287 432766 508704 432800
rect 508738 432766 508757 432800
rect 508287 432732 508306 432766
rect 508340 432750 508757 432766
rect 508340 432732 508453 432750
rect 508287 432716 508453 432732
rect 508487 432716 508554 432750
rect 508588 432716 508757 432750
rect 508287 432710 508757 432716
rect 508287 432676 508704 432710
rect 508738 432676 508757 432710
rect 508287 432642 508306 432676
rect 508340 432660 508757 432676
rect 508340 432642 508453 432660
rect 508287 432626 508453 432642
rect 508487 432626 508554 432660
rect 508588 432626 508757 432660
rect 508287 432620 508757 432626
rect 508287 432586 508704 432620
rect 508738 432586 508757 432620
rect 508287 432552 508306 432586
rect 508340 432570 508757 432586
rect 508340 432552 508453 432570
rect 508287 432536 508453 432552
rect 508487 432536 508554 432570
rect 508588 432536 508757 432570
rect 508287 432530 508757 432536
rect 508287 432496 508704 432530
rect 508738 432496 508757 432530
rect 508287 432462 508306 432496
rect 508340 432480 508757 432496
rect 508340 432462 508453 432480
rect 508287 432446 508453 432462
rect 508487 432446 508554 432480
rect 508588 432446 508757 432480
rect 508287 432440 508757 432446
rect 508287 432406 508704 432440
rect 508738 432406 508757 432440
rect 508287 432372 508306 432406
rect 508340 432390 508757 432406
rect 508340 432372 508453 432390
rect 508287 432356 508453 432372
rect 508487 432356 508554 432390
rect 508588 432356 508757 432390
rect 508287 432350 508757 432356
rect 506999 432282 507018 432316
rect 507052 432300 507469 432316
rect 507052 432282 507165 432300
rect 506999 432277 507165 432282
rect 506012 432266 507165 432277
rect 507199 432266 507266 432300
rect 507300 432277 507469 432300
rect 508287 432316 508704 432350
rect 508738 432316 508757 432350
rect 508819 432972 509513 433033
rect 508819 432938 508880 432972
rect 508914 432960 508970 432972
rect 509004 432960 509060 432972
rect 509094 432960 509150 432972
rect 508926 432938 508970 432960
rect 509026 432938 509060 432960
rect 509126 432938 509150 432960
rect 509184 432960 509240 432972
rect 509184 432938 509192 432960
rect 508819 432926 508892 432938
rect 508926 432926 508992 432938
rect 509026 432926 509092 432938
rect 509126 432926 509192 432938
rect 509226 432938 509240 432960
rect 509274 432960 509330 432972
rect 509274 432938 509292 432960
rect 509226 432926 509292 432938
rect 509326 432938 509330 432960
rect 509364 432960 509420 432972
rect 509364 432938 509392 432960
rect 509454 432938 509513 432972
rect 509326 432926 509392 432938
rect 509426 432926 509513 432938
rect 508819 432882 509513 432926
rect 508819 432848 508880 432882
rect 508914 432860 508970 432882
rect 509004 432860 509060 432882
rect 509094 432860 509150 432882
rect 508926 432848 508970 432860
rect 509026 432848 509060 432860
rect 509126 432848 509150 432860
rect 509184 432860 509240 432882
rect 509184 432848 509192 432860
rect 508819 432826 508892 432848
rect 508926 432826 508992 432848
rect 509026 432826 509092 432848
rect 509126 432826 509192 432848
rect 509226 432848 509240 432860
rect 509274 432860 509330 432882
rect 509274 432848 509292 432860
rect 509226 432826 509292 432848
rect 509326 432848 509330 432860
rect 509364 432860 509420 432882
rect 509364 432848 509392 432860
rect 509454 432848 509513 432882
rect 509326 432826 509392 432848
rect 509426 432826 509513 432848
rect 508819 432792 509513 432826
rect 508819 432758 508880 432792
rect 508914 432760 508970 432792
rect 509004 432760 509060 432792
rect 509094 432760 509150 432792
rect 508926 432758 508970 432760
rect 509026 432758 509060 432760
rect 509126 432758 509150 432760
rect 509184 432760 509240 432792
rect 509184 432758 509192 432760
rect 508819 432726 508892 432758
rect 508926 432726 508992 432758
rect 509026 432726 509092 432758
rect 509126 432726 509192 432758
rect 509226 432758 509240 432760
rect 509274 432760 509330 432792
rect 509274 432758 509292 432760
rect 509226 432726 509292 432758
rect 509326 432758 509330 432760
rect 509364 432760 509420 432792
rect 509364 432758 509392 432760
rect 509454 432758 509513 432792
rect 509326 432726 509392 432758
rect 509426 432726 509513 432758
rect 508819 432702 509513 432726
rect 508819 432668 508880 432702
rect 508914 432668 508970 432702
rect 509004 432668 509060 432702
rect 509094 432668 509150 432702
rect 509184 432668 509240 432702
rect 509274 432668 509330 432702
rect 509364 432668 509420 432702
rect 509454 432668 509513 432702
rect 508819 432660 509513 432668
rect 508819 432626 508892 432660
rect 508926 432626 508992 432660
rect 509026 432626 509092 432660
rect 509126 432626 509192 432660
rect 509226 432626 509292 432660
rect 509326 432626 509392 432660
rect 509426 432626 509513 432660
rect 508819 432612 509513 432626
rect 508819 432578 508880 432612
rect 508914 432578 508970 432612
rect 509004 432578 509060 432612
rect 509094 432578 509150 432612
rect 509184 432578 509240 432612
rect 509274 432578 509330 432612
rect 509364 432578 509420 432612
rect 509454 432578 509513 432612
rect 508819 432560 509513 432578
rect 508819 432526 508892 432560
rect 508926 432526 508992 432560
rect 509026 432526 509092 432560
rect 509126 432526 509192 432560
rect 509226 432526 509292 432560
rect 509326 432526 509392 432560
rect 509426 432526 509513 432560
rect 508819 432522 509513 432526
rect 508819 432488 508880 432522
rect 508914 432488 508970 432522
rect 509004 432488 509060 432522
rect 509094 432488 509150 432522
rect 509184 432488 509240 432522
rect 509274 432488 509330 432522
rect 509364 432488 509420 432522
rect 509454 432488 509513 432522
rect 508819 432460 509513 432488
rect 508819 432432 508892 432460
rect 508926 432432 508992 432460
rect 509026 432432 509092 432460
rect 509126 432432 509192 432460
rect 508819 432398 508880 432432
rect 508926 432426 508970 432432
rect 509026 432426 509060 432432
rect 509126 432426 509150 432432
rect 508914 432398 508970 432426
rect 509004 432398 509060 432426
rect 509094 432398 509150 432426
rect 509184 432426 509192 432432
rect 509226 432432 509292 432460
rect 509226 432426 509240 432432
rect 509184 432398 509240 432426
rect 509274 432426 509292 432432
rect 509326 432432 509392 432460
rect 509426 432432 509513 432460
rect 509326 432426 509330 432432
rect 509274 432398 509330 432426
rect 509364 432426 509392 432432
rect 509364 432398 509420 432426
rect 509454 432398 509513 432432
rect 508819 432339 509513 432398
rect 509575 433002 509594 433036
rect 509628 433020 510045 433036
rect 510863 433076 511029 433095
rect 511063 433076 511130 433110
rect 511164 433095 512317 433110
rect 511164 433076 511333 433095
rect 510863 433070 511333 433076
rect 510863 433036 511280 433070
rect 511314 433036 511333 433070
rect 509628 433002 509741 433020
rect 509575 432986 509741 433002
rect 509775 432986 509842 433020
rect 509876 432986 510045 433020
rect 509575 432980 510045 432986
rect 509575 432946 509992 432980
rect 510026 432946 510045 432980
rect 509575 432912 509594 432946
rect 509628 432930 510045 432946
rect 509628 432912 509741 432930
rect 509575 432896 509741 432912
rect 509775 432896 509842 432930
rect 509876 432896 510045 432930
rect 509575 432890 510045 432896
rect 509575 432856 509992 432890
rect 510026 432856 510045 432890
rect 509575 432822 509594 432856
rect 509628 432840 510045 432856
rect 509628 432822 509741 432840
rect 509575 432806 509741 432822
rect 509775 432806 509842 432840
rect 509876 432806 510045 432840
rect 509575 432800 510045 432806
rect 509575 432766 509992 432800
rect 510026 432766 510045 432800
rect 509575 432732 509594 432766
rect 509628 432750 510045 432766
rect 509628 432732 509741 432750
rect 509575 432716 509741 432732
rect 509775 432716 509842 432750
rect 509876 432716 510045 432750
rect 509575 432710 510045 432716
rect 509575 432676 509992 432710
rect 510026 432676 510045 432710
rect 509575 432642 509594 432676
rect 509628 432660 510045 432676
rect 509628 432642 509741 432660
rect 509575 432626 509741 432642
rect 509775 432626 509842 432660
rect 509876 432626 510045 432660
rect 509575 432620 510045 432626
rect 509575 432586 509992 432620
rect 510026 432586 510045 432620
rect 509575 432552 509594 432586
rect 509628 432570 510045 432586
rect 509628 432552 509741 432570
rect 509575 432536 509741 432552
rect 509775 432536 509842 432570
rect 509876 432536 510045 432570
rect 509575 432530 510045 432536
rect 509575 432496 509992 432530
rect 510026 432496 510045 432530
rect 509575 432462 509594 432496
rect 509628 432480 510045 432496
rect 509628 432462 509741 432480
rect 509575 432446 509741 432462
rect 509775 432446 509842 432480
rect 509876 432446 510045 432480
rect 509575 432440 510045 432446
rect 509575 432406 509992 432440
rect 510026 432406 510045 432440
rect 509575 432372 509594 432406
rect 509628 432390 510045 432406
rect 509628 432372 509741 432390
rect 509575 432356 509741 432372
rect 509775 432356 509842 432390
rect 509876 432356 510045 432390
rect 509575 432350 510045 432356
rect 508287 432282 508306 432316
rect 508340 432300 508757 432316
rect 508340 432282 508453 432300
rect 508287 432277 508453 432282
rect 507300 432266 508453 432277
rect 508487 432266 508554 432300
rect 508588 432277 508757 432300
rect 509575 432316 509992 432350
rect 510026 432316 510045 432350
rect 510107 432972 510801 433033
rect 510107 432938 510168 432972
rect 510202 432960 510258 432972
rect 510292 432960 510348 432972
rect 510382 432960 510438 432972
rect 510214 432938 510258 432960
rect 510314 432938 510348 432960
rect 510414 432938 510438 432960
rect 510472 432960 510528 432972
rect 510472 432938 510480 432960
rect 510107 432926 510180 432938
rect 510214 432926 510280 432938
rect 510314 432926 510380 432938
rect 510414 432926 510480 432938
rect 510514 432938 510528 432960
rect 510562 432960 510618 432972
rect 510562 432938 510580 432960
rect 510514 432926 510580 432938
rect 510614 432938 510618 432960
rect 510652 432960 510708 432972
rect 510652 432938 510680 432960
rect 510742 432938 510801 432972
rect 510614 432926 510680 432938
rect 510714 432926 510801 432938
rect 510107 432882 510801 432926
rect 510107 432848 510168 432882
rect 510202 432860 510258 432882
rect 510292 432860 510348 432882
rect 510382 432860 510438 432882
rect 510214 432848 510258 432860
rect 510314 432848 510348 432860
rect 510414 432848 510438 432860
rect 510472 432860 510528 432882
rect 510472 432848 510480 432860
rect 510107 432826 510180 432848
rect 510214 432826 510280 432848
rect 510314 432826 510380 432848
rect 510414 432826 510480 432848
rect 510514 432848 510528 432860
rect 510562 432860 510618 432882
rect 510562 432848 510580 432860
rect 510514 432826 510580 432848
rect 510614 432848 510618 432860
rect 510652 432860 510708 432882
rect 510652 432848 510680 432860
rect 510742 432848 510801 432882
rect 510614 432826 510680 432848
rect 510714 432826 510801 432848
rect 510107 432792 510801 432826
rect 510107 432758 510168 432792
rect 510202 432760 510258 432792
rect 510292 432760 510348 432792
rect 510382 432760 510438 432792
rect 510214 432758 510258 432760
rect 510314 432758 510348 432760
rect 510414 432758 510438 432760
rect 510472 432760 510528 432792
rect 510472 432758 510480 432760
rect 510107 432726 510180 432758
rect 510214 432726 510280 432758
rect 510314 432726 510380 432758
rect 510414 432726 510480 432758
rect 510514 432758 510528 432760
rect 510562 432760 510618 432792
rect 510562 432758 510580 432760
rect 510514 432726 510580 432758
rect 510614 432758 510618 432760
rect 510652 432760 510708 432792
rect 510652 432758 510680 432760
rect 510742 432758 510801 432792
rect 510614 432726 510680 432758
rect 510714 432726 510801 432758
rect 510107 432702 510801 432726
rect 510107 432668 510168 432702
rect 510202 432668 510258 432702
rect 510292 432668 510348 432702
rect 510382 432668 510438 432702
rect 510472 432668 510528 432702
rect 510562 432668 510618 432702
rect 510652 432668 510708 432702
rect 510742 432668 510801 432702
rect 510107 432660 510801 432668
rect 510107 432626 510180 432660
rect 510214 432626 510280 432660
rect 510314 432626 510380 432660
rect 510414 432626 510480 432660
rect 510514 432626 510580 432660
rect 510614 432626 510680 432660
rect 510714 432626 510801 432660
rect 510107 432612 510801 432626
rect 510107 432578 510168 432612
rect 510202 432578 510258 432612
rect 510292 432578 510348 432612
rect 510382 432578 510438 432612
rect 510472 432578 510528 432612
rect 510562 432578 510618 432612
rect 510652 432578 510708 432612
rect 510742 432578 510801 432612
rect 510107 432560 510801 432578
rect 510107 432526 510180 432560
rect 510214 432526 510280 432560
rect 510314 432526 510380 432560
rect 510414 432526 510480 432560
rect 510514 432526 510580 432560
rect 510614 432526 510680 432560
rect 510714 432526 510801 432560
rect 510107 432522 510801 432526
rect 510107 432488 510168 432522
rect 510202 432488 510258 432522
rect 510292 432488 510348 432522
rect 510382 432488 510438 432522
rect 510472 432488 510528 432522
rect 510562 432488 510618 432522
rect 510652 432488 510708 432522
rect 510742 432488 510801 432522
rect 510107 432460 510801 432488
rect 510107 432432 510180 432460
rect 510214 432432 510280 432460
rect 510314 432432 510380 432460
rect 510414 432432 510480 432460
rect 510107 432398 510168 432432
rect 510214 432426 510258 432432
rect 510314 432426 510348 432432
rect 510414 432426 510438 432432
rect 510202 432398 510258 432426
rect 510292 432398 510348 432426
rect 510382 432398 510438 432426
rect 510472 432426 510480 432432
rect 510514 432432 510580 432460
rect 510514 432426 510528 432432
rect 510472 432398 510528 432426
rect 510562 432426 510580 432432
rect 510614 432432 510680 432460
rect 510714 432432 510801 432460
rect 510614 432426 510618 432432
rect 510562 432398 510618 432426
rect 510652 432426 510680 432432
rect 510652 432398 510708 432426
rect 510742 432398 510801 432432
rect 510107 432339 510801 432398
rect 510863 433002 510882 433036
rect 510916 433020 511333 433036
rect 512151 433076 512317 433095
rect 512351 433076 512418 433110
rect 512452 433095 513605 433110
rect 512452 433076 512621 433095
rect 512151 433070 512621 433076
rect 512151 433036 512568 433070
rect 512602 433036 512621 433070
rect 510916 433002 511029 433020
rect 510863 432986 511029 433002
rect 511063 432986 511130 433020
rect 511164 432986 511333 433020
rect 510863 432980 511333 432986
rect 510863 432946 511280 432980
rect 511314 432946 511333 432980
rect 510863 432912 510882 432946
rect 510916 432930 511333 432946
rect 510916 432912 511029 432930
rect 510863 432896 511029 432912
rect 511063 432896 511130 432930
rect 511164 432896 511333 432930
rect 510863 432890 511333 432896
rect 510863 432856 511280 432890
rect 511314 432856 511333 432890
rect 510863 432822 510882 432856
rect 510916 432840 511333 432856
rect 510916 432822 511029 432840
rect 510863 432806 511029 432822
rect 511063 432806 511130 432840
rect 511164 432806 511333 432840
rect 510863 432800 511333 432806
rect 510863 432766 511280 432800
rect 511314 432766 511333 432800
rect 510863 432732 510882 432766
rect 510916 432750 511333 432766
rect 510916 432732 511029 432750
rect 510863 432716 511029 432732
rect 511063 432716 511130 432750
rect 511164 432716 511333 432750
rect 510863 432710 511333 432716
rect 510863 432676 511280 432710
rect 511314 432676 511333 432710
rect 510863 432642 510882 432676
rect 510916 432660 511333 432676
rect 510916 432642 511029 432660
rect 510863 432626 511029 432642
rect 511063 432626 511130 432660
rect 511164 432626 511333 432660
rect 510863 432620 511333 432626
rect 510863 432586 511280 432620
rect 511314 432586 511333 432620
rect 510863 432552 510882 432586
rect 510916 432570 511333 432586
rect 510916 432552 511029 432570
rect 510863 432536 511029 432552
rect 511063 432536 511130 432570
rect 511164 432536 511333 432570
rect 510863 432530 511333 432536
rect 510863 432496 511280 432530
rect 511314 432496 511333 432530
rect 510863 432462 510882 432496
rect 510916 432480 511333 432496
rect 510916 432462 511029 432480
rect 510863 432446 511029 432462
rect 511063 432446 511130 432480
rect 511164 432446 511333 432480
rect 510863 432440 511333 432446
rect 510863 432406 511280 432440
rect 511314 432406 511333 432440
rect 510863 432372 510882 432406
rect 510916 432390 511333 432406
rect 510916 432372 511029 432390
rect 510863 432356 511029 432372
rect 511063 432356 511130 432390
rect 511164 432356 511333 432390
rect 510863 432350 511333 432356
rect 509575 432282 509594 432316
rect 509628 432300 510045 432316
rect 509628 432282 509741 432300
rect 509575 432277 509741 432282
rect 508588 432266 509741 432277
rect 509775 432266 509842 432300
rect 509876 432277 510045 432300
rect 510863 432316 511280 432350
rect 511314 432316 511333 432350
rect 511395 432972 512089 433033
rect 511395 432938 511456 432972
rect 511490 432960 511546 432972
rect 511580 432960 511636 432972
rect 511670 432960 511726 432972
rect 511502 432938 511546 432960
rect 511602 432938 511636 432960
rect 511702 432938 511726 432960
rect 511760 432960 511816 432972
rect 511760 432938 511768 432960
rect 511395 432926 511468 432938
rect 511502 432926 511568 432938
rect 511602 432926 511668 432938
rect 511702 432926 511768 432938
rect 511802 432938 511816 432960
rect 511850 432960 511906 432972
rect 511850 432938 511868 432960
rect 511802 432926 511868 432938
rect 511902 432938 511906 432960
rect 511940 432960 511996 432972
rect 511940 432938 511968 432960
rect 512030 432938 512089 432972
rect 511902 432926 511968 432938
rect 512002 432926 512089 432938
rect 511395 432882 512089 432926
rect 511395 432848 511456 432882
rect 511490 432860 511546 432882
rect 511580 432860 511636 432882
rect 511670 432860 511726 432882
rect 511502 432848 511546 432860
rect 511602 432848 511636 432860
rect 511702 432848 511726 432860
rect 511760 432860 511816 432882
rect 511760 432848 511768 432860
rect 511395 432826 511468 432848
rect 511502 432826 511568 432848
rect 511602 432826 511668 432848
rect 511702 432826 511768 432848
rect 511802 432848 511816 432860
rect 511850 432860 511906 432882
rect 511850 432848 511868 432860
rect 511802 432826 511868 432848
rect 511902 432848 511906 432860
rect 511940 432860 511996 432882
rect 511940 432848 511968 432860
rect 512030 432848 512089 432882
rect 511902 432826 511968 432848
rect 512002 432826 512089 432848
rect 511395 432792 512089 432826
rect 511395 432758 511456 432792
rect 511490 432760 511546 432792
rect 511580 432760 511636 432792
rect 511670 432760 511726 432792
rect 511502 432758 511546 432760
rect 511602 432758 511636 432760
rect 511702 432758 511726 432760
rect 511760 432760 511816 432792
rect 511760 432758 511768 432760
rect 511395 432726 511468 432758
rect 511502 432726 511568 432758
rect 511602 432726 511668 432758
rect 511702 432726 511768 432758
rect 511802 432758 511816 432760
rect 511850 432760 511906 432792
rect 511850 432758 511868 432760
rect 511802 432726 511868 432758
rect 511902 432758 511906 432760
rect 511940 432760 511996 432792
rect 511940 432758 511968 432760
rect 512030 432758 512089 432792
rect 511902 432726 511968 432758
rect 512002 432726 512089 432758
rect 511395 432702 512089 432726
rect 511395 432668 511456 432702
rect 511490 432668 511546 432702
rect 511580 432668 511636 432702
rect 511670 432668 511726 432702
rect 511760 432668 511816 432702
rect 511850 432668 511906 432702
rect 511940 432668 511996 432702
rect 512030 432668 512089 432702
rect 511395 432660 512089 432668
rect 511395 432626 511468 432660
rect 511502 432626 511568 432660
rect 511602 432626 511668 432660
rect 511702 432626 511768 432660
rect 511802 432626 511868 432660
rect 511902 432626 511968 432660
rect 512002 432626 512089 432660
rect 511395 432612 512089 432626
rect 511395 432578 511456 432612
rect 511490 432578 511546 432612
rect 511580 432578 511636 432612
rect 511670 432578 511726 432612
rect 511760 432578 511816 432612
rect 511850 432578 511906 432612
rect 511940 432578 511996 432612
rect 512030 432578 512089 432612
rect 511395 432560 512089 432578
rect 511395 432526 511468 432560
rect 511502 432526 511568 432560
rect 511602 432526 511668 432560
rect 511702 432526 511768 432560
rect 511802 432526 511868 432560
rect 511902 432526 511968 432560
rect 512002 432526 512089 432560
rect 511395 432522 512089 432526
rect 511395 432488 511456 432522
rect 511490 432488 511546 432522
rect 511580 432488 511636 432522
rect 511670 432488 511726 432522
rect 511760 432488 511816 432522
rect 511850 432488 511906 432522
rect 511940 432488 511996 432522
rect 512030 432488 512089 432522
rect 511395 432460 512089 432488
rect 511395 432432 511468 432460
rect 511502 432432 511568 432460
rect 511602 432432 511668 432460
rect 511702 432432 511768 432460
rect 511395 432398 511456 432432
rect 511502 432426 511546 432432
rect 511602 432426 511636 432432
rect 511702 432426 511726 432432
rect 511490 432398 511546 432426
rect 511580 432398 511636 432426
rect 511670 432398 511726 432426
rect 511760 432426 511768 432432
rect 511802 432432 511868 432460
rect 511802 432426 511816 432432
rect 511760 432398 511816 432426
rect 511850 432426 511868 432432
rect 511902 432432 511968 432460
rect 512002 432432 512089 432460
rect 511902 432426 511906 432432
rect 511850 432398 511906 432426
rect 511940 432426 511968 432432
rect 511940 432398 511996 432426
rect 512030 432398 512089 432432
rect 511395 432339 512089 432398
rect 512151 433002 512170 433036
rect 512204 433020 512621 433036
rect 513439 433076 513605 433095
rect 513639 433076 513674 433110
rect 513439 433036 513674 433076
rect 512204 433002 512317 433020
rect 512151 432986 512317 433002
rect 512351 432986 512418 433020
rect 512452 432986 512621 433020
rect 512151 432980 512621 432986
rect 512151 432946 512568 432980
rect 512602 432946 512621 432980
rect 512151 432912 512170 432946
rect 512204 432930 512621 432946
rect 512204 432912 512317 432930
rect 512151 432896 512317 432912
rect 512351 432896 512418 432930
rect 512452 432896 512621 432930
rect 512151 432890 512621 432896
rect 512151 432856 512568 432890
rect 512602 432856 512621 432890
rect 512151 432822 512170 432856
rect 512204 432840 512621 432856
rect 512204 432822 512317 432840
rect 512151 432806 512317 432822
rect 512351 432806 512418 432840
rect 512452 432806 512621 432840
rect 512151 432800 512621 432806
rect 512151 432766 512568 432800
rect 512602 432766 512621 432800
rect 512151 432732 512170 432766
rect 512204 432750 512621 432766
rect 512204 432732 512317 432750
rect 512151 432716 512317 432732
rect 512351 432716 512418 432750
rect 512452 432716 512621 432750
rect 512151 432710 512621 432716
rect 512151 432676 512568 432710
rect 512602 432676 512621 432710
rect 512151 432642 512170 432676
rect 512204 432660 512621 432676
rect 512204 432642 512317 432660
rect 512151 432626 512317 432642
rect 512351 432626 512418 432660
rect 512452 432626 512621 432660
rect 512151 432620 512621 432626
rect 512151 432586 512568 432620
rect 512602 432586 512621 432620
rect 512151 432552 512170 432586
rect 512204 432570 512621 432586
rect 512204 432552 512317 432570
rect 512151 432536 512317 432552
rect 512351 432536 512418 432570
rect 512452 432536 512621 432570
rect 512151 432530 512621 432536
rect 512151 432496 512568 432530
rect 512602 432496 512621 432530
rect 512151 432462 512170 432496
rect 512204 432480 512621 432496
rect 512204 432462 512317 432480
rect 512151 432446 512317 432462
rect 512351 432446 512418 432480
rect 512452 432446 512621 432480
rect 512151 432440 512621 432446
rect 512151 432406 512568 432440
rect 512602 432406 512621 432440
rect 512151 432372 512170 432406
rect 512204 432390 512621 432406
rect 512204 432372 512317 432390
rect 512151 432356 512317 432372
rect 512351 432356 512418 432390
rect 512452 432356 512621 432390
rect 512151 432350 512621 432356
rect 510863 432282 510882 432316
rect 510916 432300 511333 432316
rect 510916 432282 511029 432300
rect 510863 432277 511029 432282
rect 509876 432266 511029 432277
rect 511063 432266 511130 432300
rect 511164 432277 511333 432300
rect 512151 432316 512568 432350
rect 512602 432316 512621 432350
rect 512683 432972 513377 433033
rect 512683 432938 512744 432972
rect 512778 432960 512834 432972
rect 512868 432960 512924 432972
rect 512958 432960 513014 432972
rect 512790 432938 512834 432960
rect 512890 432938 512924 432960
rect 512990 432938 513014 432960
rect 513048 432960 513104 432972
rect 513048 432938 513056 432960
rect 512683 432926 512756 432938
rect 512790 432926 512856 432938
rect 512890 432926 512956 432938
rect 512990 432926 513056 432938
rect 513090 432938 513104 432960
rect 513138 432960 513194 432972
rect 513138 432938 513156 432960
rect 513090 432926 513156 432938
rect 513190 432938 513194 432960
rect 513228 432960 513284 432972
rect 513228 432938 513256 432960
rect 513318 432938 513377 432972
rect 513190 432926 513256 432938
rect 513290 432926 513377 432938
rect 512683 432882 513377 432926
rect 512683 432848 512744 432882
rect 512778 432860 512834 432882
rect 512868 432860 512924 432882
rect 512958 432860 513014 432882
rect 512790 432848 512834 432860
rect 512890 432848 512924 432860
rect 512990 432848 513014 432860
rect 513048 432860 513104 432882
rect 513048 432848 513056 432860
rect 512683 432826 512756 432848
rect 512790 432826 512856 432848
rect 512890 432826 512956 432848
rect 512990 432826 513056 432848
rect 513090 432848 513104 432860
rect 513138 432860 513194 432882
rect 513138 432848 513156 432860
rect 513090 432826 513156 432848
rect 513190 432848 513194 432860
rect 513228 432860 513284 432882
rect 513228 432848 513256 432860
rect 513318 432848 513377 432882
rect 513190 432826 513256 432848
rect 513290 432826 513377 432848
rect 512683 432792 513377 432826
rect 512683 432758 512744 432792
rect 512778 432760 512834 432792
rect 512868 432760 512924 432792
rect 512958 432760 513014 432792
rect 512790 432758 512834 432760
rect 512890 432758 512924 432760
rect 512990 432758 513014 432760
rect 513048 432760 513104 432792
rect 513048 432758 513056 432760
rect 512683 432726 512756 432758
rect 512790 432726 512856 432758
rect 512890 432726 512956 432758
rect 512990 432726 513056 432758
rect 513090 432758 513104 432760
rect 513138 432760 513194 432792
rect 513138 432758 513156 432760
rect 513090 432726 513156 432758
rect 513190 432758 513194 432760
rect 513228 432760 513284 432792
rect 513228 432758 513256 432760
rect 513318 432758 513377 432792
rect 513190 432726 513256 432758
rect 513290 432726 513377 432758
rect 512683 432702 513377 432726
rect 512683 432668 512744 432702
rect 512778 432668 512834 432702
rect 512868 432668 512924 432702
rect 512958 432668 513014 432702
rect 513048 432668 513104 432702
rect 513138 432668 513194 432702
rect 513228 432668 513284 432702
rect 513318 432668 513377 432702
rect 512683 432660 513377 432668
rect 512683 432626 512756 432660
rect 512790 432626 512856 432660
rect 512890 432626 512956 432660
rect 512990 432626 513056 432660
rect 513090 432626 513156 432660
rect 513190 432626 513256 432660
rect 513290 432626 513377 432660
rect 512683 432612 513377 432626
rect 512683 432578 512744 432612
rect 512778 432578 512834 432612
rect 512868 432578 512924 432612
rect 512958 432578 513014 432612
rect 513048 432578 513104 432612
rect 513138 432578 513194 432612
rect 513228 432578 513284 432612
rect 513318 432578 513377 432612
rect 512683 432560 513377 432578
rect 512683 432526 512756 432560
rect 512790 432526 512856 432560
rect 512890 432526 512956 432560
rect 512990 432526 513056 432560
rect 513090 432526 513156 432560
rect 513190 432526 513256 432560
rect 513290 432526 513377 432560
rect 512683 432522 513377 432526
rect 512683 432488 512744 432522
rect 512778 432488 512834 432522
rect 512868 432488 512924 432522
rect 512958 432488 513014 432522
rect 513048 432488 513104 432522
rect 513138 432488 513194 432522
rect 513228 432488 513284 432522
rect 513318 432488 513377 432522
rect 512683 432460 513377 432488
rect 512683 432432 512756 432460
rect 512790 432432 512856 432460
rect 512890 432432 512956 432460
rect 512990 432432 513056 432460
rect 512683 432398 512744 432432
rect 512790 432426 512834 432432
rect 512890 432426 512924 432432
rect 512990 432426 513014 432432
rect 512778 432398 512834 432426
rect 512868 432398 512924 432426
rect 512958 432398 513014 432426
rect 513048 432426 513056 432432
rect 513090 432432 513156 432460
rect 513090 432426 513104 432432
rect 513048 432398 513104 432426
rect 513138 432426 513156 432432
rect 513190 432432 513256 432460
rect 513290 432432 513377 432460
rect 513190 432426 513194 432432
rect 513138 432398 513194 432426
rect 513228 432426 513256 432432
rect 513228 432398 513284 432426
rect 513318 432398 513377 432432
rect 512683 432339 513377 432398
rect 513439 433002 513458 433036
rect 513492 433020 513674 433036
rect 513492 433002 513605 433020
rect 513439 432986 513605 433002
rect 513639 432986 513674 433020
rect 513439 432946 513674 432986
rect 513439 432912 513458 432946
rect 513492 432930 513674 432946
rect 513492 432912 513605 432930
rect 513439 432896 513605 432912
rect 513639 432896 513674 432930
rect 513439 432856 513674 432896
rect 513439 432822 513458 432856
rect 513492 432840 513674 432856
rect 513492 432822 513605 432840
rect 513439 432806 513605 432822
rect 513639 432806 513674 432840
rect 513439 432766 513674 432806
rect 513439 432732 513458 432766
rect 513492 432750 513674 432766
rect 513492 432732 513605 432750
rect 513439 432716 513605 432732
rect 513639 432716 513674 432750
rect 513439 432676 513674 432716
rect 513439 432642 513458 432676
rect 513492 432660 513674 432676
rect 513492 432642 513605 432660
rect 513439 432626 513605 432642
rect 513639 432626 513674 432660
rect 513439 432586 513674 432626
rect 513439 432552 513458 432586
rect 513492 432570 513674 432586
rect 513492 432552 513605 432570
rect 513439 432536 513605 432552
rect 513639 432536 513674 432570
rect 513439 432496 513674 432536
rect 513439 432462 513458 432496
rect 513492 432480 513674 432496
rect 513492 432462 513605 432480
rect 513439 432446 513605 432462
rect 513639 432446 513674 432480
rect 513439 432406 513674 432446
rect 513439 432372 513458 432406
rect 513492 432390 513674 432406
rect 513492 432372 513605 432390
rect 513439 432356 513605 432372
rect 513639 432356 513674 432390
rect 512151 432282 512170 432316
rect 512204 432300 512621 432316
rect 512204 432282 512317 432300
rect 512151 432277 512317 432282
rect 511164 432266 512317 432277
rect 512351 432266 512418 432300
rect 512452 432277 512621 432300
rect 513439 432316 513674 432356
rect 513439 432282 513458 432316
rect 513492 432300 513674 432316
rect 513492 432282 513605 432300
rect 513439 432277 513605 432282
rect 512452 432266 513605 432277
rect 513639 432266 513674 432300
rect 503370 432258 513674 432266
rect 503370 432224 503646 432258
rect 503680 432224 503736 432258
rect 503770 432224 503826 432258
rect 503860 432224 503916 432258
rect 503950 432224 504006 432258
rect 504040 432224 504096 432258
rect 504130 432224 504186 432258
rect 504220 432224 504276 432258
rect 504310 432224 504366 432258
rect 504400 432224 504934 432258
rect 504968 432224 505024 432258
rect 505058 432224 505114 432258
rect 505148 432224 505204 432258
rect 505238 432224 505294 432258
rect 505328 432224 505384 432258
rect 505418 432224 505474 432258
rect 505508 432224 505564 432258
rect 505598 432224 505654 432258
rect 505688 432224 506222 432258
rect 506256 432224 506312 432258
rect 506346 432224 506402 432258
rect 506436 432224 506492 432258
rect 506526 432224 506582 432258
rect 506616 432224 506672 432258
rect 506706 432224 506762 432258
rect 506796 432224 506852 432258
rect 506886 432224 506942 432258
rect 506976 432224 507510 432258
rect 507544 432224 507600 432258
rect 507634 432224 507690 432258
rect 507724 432224 507780 432258
rect 507814 432224 507870 432258
rect 507904 432224 507960 432258
rect 507994 432224 508050 432258
rect 508084 432224 508140 432258
rect 508174 432224 508230 432258
rect 508264 432224 508798 432258
rect 508832 432224 508888 432258
rect 508922 432224 508978 432258
rect 509012 432224 509068 432258
rect 509102 432224 509158 432258
rect 509192 432224 509248 432258
rect 509282 432224 509338 432258
rect 509372 432224 509428 432258
rect 509462 432224 509518 432258
rect 509552 432224 510086 432258
rect 510120 432224 510176 432258
rect 510210 432224 510266 432258
rect 510300 432224 510356 432258
rect 510390 432224 510446 432258
rect 510480 432224 510536 432258
rect 510570 432224 510626 432258
rect 510660 432224 510716 432258
rect 510750 432224 510806 432258
rect 510840 432224 511374 432258
rect 511408 432224 511464 432258
rect 511498 432224 511554 432258
rect 511588 432224 511644 432258
rect 511678 432224 511734 432258
rect 511768 432224 511824 432258
rect 511858 432224 511914 432258
rect 511948 432224 512004 432258
rect 512038 432224 512094 432258
rect 512128 432224 512662 432258
rect 512696 432224 512752 432258
rect 512786 432224 512842 432258
rect 512876 432224 512932 432258
rect 512966 432224 513022 432258
rect 513056 432224 513112 432258
rect 513146 432224 513202 432258
rect 513236 432224 513292 432258
rect 513326 432224 513382 432258
rect 513416 432224 513674 432258
rect 503370 432210 513674 432224
rect 503370 432176 503402 432210
rect 503436 432176 504589 432210
rect 504623 432176 504690 432210
rect 504724 432176 505877 432210
rect 505911 432176 505978 432210
rect 506012 432176 507165 432210
rect 507199 432176 507266 432210
rect 507300 432176 508453 432210
rect 508487 432176 508554 432210
rect 508588 432176 509741 432210
rect 509775 432176 509842 432210
rect 509876 432176 511029 432210
rect 511063 432176 511130 432210
rect 511164 432176 512317 432210
rect 512351 432176 512418 432210
rect 512452 432176 513605 432210
rect 513639 432176 513674 432210
rect 500320 432064 500418 432068
rect 500518 432064 500642 432068
rect 500742 432064 500866 432068
rect 500966 432064 501090 432068
rect 501190 432064 501314 432068
rect 503370 432109 513674 432176
rect 503370 432075 503486 432109
rect 503520 432075 503576 432109
rect 503610 432075 503666 432109
rect 503700 432075 503756 432109
rect 503790 432075 503846 432109
rect 503880 432075 503936 432109
rect 503970 432075 504026 432109
rect 504060 432075 504116 432109
rect 504150 432075 504206 432109
rect 504240 432075 504296 432109
rect 504330 432075 504386 432109
rect 504420 432075 504476 432109
rect 504510 432075 504566 432109
rect 504600 432075 504774 432109
rect 504808 432075 504864 432109
rect 504898 432075 504954 432109
rect 504988 432075 505044 432109
rect 505078 432075 505134 432109
rect 505168 432075 505224 432109
rect 505258 432075 505314 432109
rect 505348 432075 505404 432109
rect 505438 432075 505494 432109
rect 505528 432075 505584 432109
rect 505618 432075 505674 432109
rect 505708 432075 505764 432109
rect 505798 432075 505854 432109
rect 505888 432075 506062 432109
rect 506096 432075 506152 432109
rect 506186 432075 506242 432109
rect 506276 432075 506332 432109
rect 506366 432075 506422 432109
rect 506456 432075 506512 432109
rect 506546 432075 506602 432109
rect 506636 432075 506692 432109
rect 506726 432075 506782 432109
rect 506816 432075 506872 432109
rect 506906 432075 506962 432109
rect 506996 432075 507052 432109
rect 507086 432075 507142 432109
rect 507176 432075 507350 432109
rect 507384 432075 507440 432109
rect 507474 432075 507530 432109
rect 507564 432075 507620 432109
rect 507654 432075 507710 432109
rect 507744 432075 507800 432109
rect 507834 432075 507890 432109
rect 507924 432075 507980 432109
rect 508014 432075 508070 432109
rect 508104 432075 508160 432109
rect 508194 432075 508250 432109
rect 508284 432075 508340 432109
rect 508374 432075 508430 432109
rect 508464 432075 508638 432109
rect 508672 432075 508728 432109
rect 508762 432075 508818 432109
rect 508852 432075 508908 432109
rect 508942 432075 508998 432109
rect 509032 432075 509088 432109
rect 509122 432075 509178 432109
rect 509212 432075 509268 432109
rect 509302 432075 509358 432109
rect 509392 432075 509448 432109
rect 509482 432075 509538 432109
rect 509572 432075 509628 432109
rect 509662 432075 509718 432109
rect 509752 432075 509926 432109
rect 509960 432075 510016 432109
rect 510050 432075 510106 432109
rect 510140 432075 510196 432109
rect 510230 432075 510286 432109
rect 510320 432075 510376 432109
rect 510410 432075 510466 432109
rect 510500 432075 510556 432109
rect 510590 432075 510646 432109
rect 510680 432075 510736 432109
rect 510770 432075 510826 432109
rect 510860 432075 510916 432109
rect 510950 432075 511006 432109
rect 511040 432075 511214 432109
rect 511248 432075 511304 432109
rect 511338 432075 511394 432109
rect 511428 432075 511484 432109
rect 511518 432075 511574 432109
rect 511608 432075 511664 432109
rect 511698 432075 511754 432109
rect 511788 432075 511844 432109
rect 511878 432075 511934 432109
rect 511968 432075 512024 432109
rect 512058 432075 512114 432109
rect 512148 432075 512204 432109
rect 512238 432075 512294 432109
rect 512328 432075 512502 432109
rect 512536 432075 512592 432109
rect 512626 432075 512682 432109
rect 512716 432075 512772 432109
rect 512806 432075 512862 432109
rect 512896 432075 512952 432109
rect 512986 432075 513042 432109
rect 513076 432075 513132 432109
rect 513166 432075 513222 432109
rect 513256 432075 513312 432109
rect 513346 432075 513402 432109
rect 513436 432075 513492 432109
rect 513526 432075 513582 432109
rect 513616 432075 513674 432109
rect 500320 432052 501384 432064
rect 500320 431940 501344 432052
rect 503370 432042 513674 432075
rect 500320 431840 500418 431940
rect 500518 431840 500642 431940
rect 500742 431840 500866 431940
rect 500966 431840 501090 431940
rect 501190 431840 501314 431940
rect 500320 431716 501344 431840
rect 500320 431616 500418 431716
rect 500518 431616 500642 431716
rect 500742 431616 500866 431716
rect 500966 431616 501090 431716
rect 501190 431616 501314 431716
rect 500320 431492 501344 431616
rect 500320 431392 500418 431492
rect 500518 431392 500642 431492
rect 500742 431392 500866 431492
rect 500966 431392 501090 431492
rect 501190 431392 501314 431492
rect 500320 431268 501344 431392
rect 500320 431168 500418 431268
rect 500518 431168 500642 431268
rect 500742 431168 500866 431268
rect 500966 431168 501090 431268
rect 501190 431168 501314 431268
rect 500320 431060 501344 431168
rect 500320 431044 526584 431060
rect 500320 430044 500344 431044
rect 526568 430996 526584 431044
rect 527576 430996 527592 474332
rect 528592 474332 528616 475332
rect 528592 474280 528608 474332
rect 528592 474056 528608 474180
rect 528592 473832 528608 473956
rect 528592 473608 528608 473732
rect 528592 473384 528608 473508
rect 528592 473160 528608 473284
rect 528592 472936 528608 473060
rect 528592 472712 528608 472836
rect 528592 472488 528608 472612
rect 528592 472264 528608 472388
rect 528592 472040 528608 472164
rect 528592 471816 528608 471940
rect 528592 471592 528608 471716
rect 528592 471368 528608 471492
rect 528592 471144 528608 471268
rect 528592 470920 528608 471044
rect 528592 470696 528608 470820
rect 528592 470472 528608 470596
rect 528592 470248 528608 470372
rect 528592 470024 528608 470148
rect 528592 469800 528608 469924
rect 528592 469576 528608 469700
rect 528592 469352 528608 469476
rect 528592 469128 528608 469252
rect 528592 468904 528608 469028
rect 528592 468680 528608 468804
rect 528592 468456 528608 468580
rect 528592 468232 528608 468356
rect 528592 468008 528608 468132
rect 528592 467784 528608 467908
rect 528592 463810 528608 467684
rect 528592 463586 528608 463710
rect 528592 463362 528608 463486
rect 528592 463138 528608 463262
rect 528592 462914 528608 463038
rect 528592 462690 528608 462814
rect 528592 462466 528608 462590
rect 528592 462242 528608 462366
rect 528592 462018 528608 462142
rect 528592 461794 528608 461918
rect 528592 461570 528608 461694
rect 528592 461346 528608 461470
rect 528592 461122 528608 461246
rect 528592 460898 528608 461022
rect 528592 460674 528608 460798
rect 528592 460450 528608 460574
rect 528592 460226 528608 460350
rect 528592 460002 528608 460126
rect 528592 459778 528608 459902
rect 528592 459554 528608 459678
rect 528592 459330 528608 459454
rect 528592 459106 528608 459230
rect 528592 458882 528608 459006
rect 528592 458658 528608 458782
rect 528592 458434 528608 458558
rect 528592 458210 528608 458334
rect 528592 457986 528608 458110
rect 528592 457762 528608 457886
rect 528592 457538 528608 457662
rect 528592 457314 528608 457438
rect 528592 437540 528608 457214
rect 562156 455115 562190 455212
rect 567544 455115 567578 455212
rect 562270 455088 562304 455104
rect 562270 454096 562304 454112
rect 562528 455088 562562 455104
rect 562528 454053 562562 454112
rect 562786 455088 562820 455104
rect 562786 454096 562820 454112
rect 563044 455088 563078 455104
rect 563044 454053 563078 454112
rect 563302 455088 563336 455104
rect 563302 454096 563336 454112
rect 563560 455088 563594 455104
rect 563560 454053 563594 454112
rect 563818 455088 563852 455104
rect 563818 454096 563852 454112
rect 564076 455088 564110 455104
rect 564076 454053 564110 454112
rect 564334 455088 564368 455104
rect 564334 454096 564368 454112
rect 564592 455088 564626 455104
rect 564592 454053 564626 454112
rect 564850 455088 564884 455104
rect 564850 454096 564884 454112
rect 565108 455088 565142 455104
rect 565108 454053 565142 454112
rect 565366 455088 565400 455104
rect 565366 454096 565400 454112
rect 565624 455088 565658 455104
rect 565624 454053 565658 454112
rect 565882 455088 565916 455104
rect 565882 454096 565916 454112
rect 566140 455088 566174 455104
rect 566140 454053 566174 454112
rect 566398 455088 566432 455104
rect 566398 454096 566432 454112
rect 566656 455088 566690 455104
rect 566656 454053 566690 454112
rect 566914 455088 566948 455104
rect 566914 454096 566948 454112
rect 567172 455088 567206 455104
rect 567172 454053 567206 454112
rect 567430 455088 567464 455104
rect 567430 454096 567464 454112
rect 562270 454019 562332 454053
rect 562500 454019 562590 454053
rect 562758 454019 562848 454053
rect 563016 454019 563106 454053
rect 563274 454019 563364 454053
rect 563532 454019 563622 454053
rect 563790 454019 563880 454053
rect 564048 454019 564138 454053
rect 564306 454019 564396 454053
rect 564564 454019 564654 454053
rect 564822 454019 564912 454053
rect 565080 454019 565170 454053
rect 565338 454019 565428 454053
rect 565596 454019 565686 454053
rect 565854 454019 565944 454053
rect 566112 454019 566202 454053
rect 566370 454019 566460 454053
rect 566628 454019 566718 454053
rect 566886 454019 566976 454053
rect 567144 454019 567234 454053
rect 567402 454019 567464 454053
rect 562156 453950 562190 454013
rect 567544 453950 567578 454013
rect 572316 455150 572350 455246
rect 577704 455150 577738 455246
rect 572430 455122 572464 455138
rect 572430 454130 572464 454146
rect 572688 455122 572722 455138
rect 572688 454096 572722 454146
rect 572946 455122 572980 455138
rect 572946 454130 572980 454146
rect 573204 455122 573238 455138
rect 573204 454096 573238 454146
rect 573462 455122 573496 455138
rect 573462 454130 573496 454146
rect 573720 455122 573754 455138
rect 573720 454096 573754 454146
rect 573978 455122 574012 455138
rect 573978 454130 574012 454146
rect 574236 455122 574270 455138
rect 574236 454096 574270 454146
rect 574494 455122 574528 455138
rect 574494 454130 574528 454146
rect 574752 455122 574786 455138
rect 574752 454096 574786 454146
rect 575010 455122 575044 455138
rect 575010 454130 575044 454146
rect 575268 455122 575302 455138
rect 575268 454096 575302 454146
rect 575526 455122 575560 455138
rect 575526 454130 575560 454146
rect 575784 455122 575818 455138
rect 575784 454096 575818 454146
rect 576042 455122 576076 455138
rect 576042 454130 576076 454146
rect 576300 455122 576334 455138
rect 576300 454096 576334 454146
rect 576558 455122 576592 455138
rect 576558 454130 576592 454146
rect 576816 455122 576850 455138
rect 576816 454096 576850 454146
rect 577074 455122 577108 455138
rect 577074 454130 577108 454146
rect 577332 455122 577366 455138
rect 577332 454096 577366 454146
rect 577590 455122 577624 455138
rect 577590 454130 577624 454146
rect 572429 454062 572492 454096
rect 572660 454062 572750 454096
rect 572918 454062 573008 454096
rect 573176 454062 573266 454096
rect 573434 454062 573524 454096
rect 573692 454062 573782 454096
rect 573950 454062 574040 454096
rect 574208 454062 574298 454096
rect 574466 454062 574556 454096
rect 574724 454062 574814 454096
rect 574982 454062 575072 454096
rect 575240 454062 575330 454096
rect 575498 454062 575588 454096
rect 575756 454062 575846 454096
rect 576014 454062 576104 454096
rect 576272 454062 576362 454096
rect 576530 454062 576620 454096
rect 576788 454062 576878 454096
rect 577046 454062 577136 454096
rect 577304 454062 577394 454096
rect 577562 454062 577626 454096
rect 572316 453994 572350 454056
rect 577704 453994 577738 454056
rect 572316 453960 572412 453994
rect 577642 453960 577738 453994
rect 562156 453916 562252 453950
rect 567482 453916 567578 453950
rect 528592 437316 528608 437440
rect 528592 437092 528608 437216
rect 528592 436868 528608 436992
rect 528592 436644 528608 436768
rect 528592 436420 528608 436544
rect 528592 436196 528608 436320
rect 528592 435972 528608 436096
rect 528592 435748 528608 435872
rect 528592 435524 528608 435648
rect 528592 435300 528608 435424
rect 528592 435076 528608 435200
rect 528592 434852 528608 434976
rect 528592 434628 528608 434752
rect 528592 434404 528608 434528
rect 528592 434180 528608 434304
rect 528592 433956 528608 434080
rect 528592 433732 528608 433856
rect 528592 433508 528608 433632
rect 528592 433284 528608 433408
rect 528592 433060 528608 433184
rect 528592 432836 528608 432960
rect 528592 432612 528608 432736
rect 528592 432388 528608 432512
rect 528592 432164 528608 432288
rect 528592 431940 528608 432064
rect 528592 431716 528608 431840
rect 528592 431492 528608 431616
rect 528592 431268 528608 431392
rect 528592 431044 528608 431168
rect 526568 430044 527592 430996
rect 500320 430030 503920 430044
rect 504020 430030 504144 430044
rect 504244 430030 504368 430044
rect 504468 430030 504592 430044
rect 504692 430030 504816 430044
rect 504916 430030 505040 430044
rect 505140 430030 505264 430044
rect 505364 430030 505488 430044
rect 505588 430030 505712 430044
rect 505812 430030 505936 430044
rect 506036 430030 506160 430044
rect 506260 430030 506384 430044
rect 506484 430030 506608 430044
rect 506708 430030 506832 430044
rect 506932 430030 507056 430044
rect 507156 430030 507280 430044
rect 507380 430030 507504 430044
rect 507604 430030 507728 430044
rect 507828 430030 507952 430044
rect 508052 430030 508176 430044
rect 508276 430030 508400 430044
rect 508500 430030 508624 430044
rect 508724 430030 508848 430044
rect 508948 430030 509072 430044
rect 509172 430030 509296 430044
rect 509396 430030 509520 430044
rect 509620 430030 509744 430044
rect 509844 430030 509968 430044
rect 510068 430030 510192 430044
rect 510292 430030 510416 430044
rect 510516 430030 517320 430044
rect 517420 430030 517544 430044
rect 517644 430030 517768 430044
rect 517868 430030 517992 430044
rect 518092 430030 518216 430044
rect 518316 430030 518440 430044
rect 518540 430030 518664 430044
rect 518764 430030 518888 430044
rect 518988 430030 519112 430044
rect 519212 430030 519336 430044
rect 519436 430030 519560 430044
rect 519660 430030 519784 430044
rect 519884 430030 520008 430044
rect 520108 430030 520232 430044
rect 520332 430030 520456 430044
rect 520556 430030 520680 430044
rect 520780 430030 520904 430044
rect 521004 430030 521128 430044
rect 521228 430030 521352 430044
rect 521452 430030 521576 430044
rect 521676 430030 521800 430044
rect 521900 430030 522024 430044
rect 522124 430030 522248 430044
rect 522348 430030 522472 430044
rect 522572 430030 522696 430044
rect 522796 430030 522920 430044
rect 523020 430030 523144 430044
rect 523244 430030 523368 430044
rect 523468 430030 523592 430044
rect 523692 430030 523816 430044
rect 523916 430030 527592 430044
rect 500320 430020 527592 430030
rect 528592 430020 528616 430944
rect 500320 429996 528616 430020
<< viali >>
rect 562190 495480 562252 495514
rect 562252 495480 567482 495514
rect 567482 495480 567544 495514
rect 562156 494375 562190 495357
rect 562270 494414 562304 495390
rect 562528 494414 562562 495390
rect 562786 494414 562820 495390
rect 563044 494414 563078 495390
rect 563302 494414 563336 495390
rect 563560 494414 563594 495390
rect 563818 494414 563852 495390
rect 564076 494414 564110 495390
rect 564334 494414 564368 495390
rect 564592 494414 564626 495390
rect 564850 494414 564884 495390
rect 565108 494414 565142 495390
rect 565366 494414 565400 495390
rect 565624 494414 565658 495390
rect 565882 494414 565916 495390
rect 566140 494414 566174 495390
rect 566398 494414 566432 495390
rect 566656 494414 566690 495390
rect 566914 494414 566948 495390
rect 567172 494414 567206 495390
rect 567430 494414 567464 495390
rect 567544 494375 567578 495357
rect 562374 494321 562458 494355
rect 562632 494321 562716 494355
rect 562890 494321 562974 494355
rect 563148 494321 563232 494355
rect 563406 494321 563490 494355
rect 563664 494321 563748 494355
rect 563922 494321 564006 494355
rect 564180 494321 564264 494355
rect 564438 494321 564522 494355
rect 564696 494321 564780 494355
rect 564954 494321 565038 494355
rect 565212 494321 565296 494355
rect 565470 494321 565554 494355
rect 565728 494321 565812 494355
rect 565986 494321 566070 494355
rect 566244 494321 566328 494355
rect 566502 494321 566586 494355
rect 566760 494321 566844 494355
rect 567018 494321 567102 494355
rect 567276 494321 567360 494355
rect 572350 495514 572412 495548
rect 572412 495514 577642 495548
rect 577642 495514 577704 495548
rect 572316 494418 572350 495392
rect 572430 494448 572464 495424
rect 572688 494448 572722 495424
rect 572946 494448 572980 495424
rect 573204 494448 573238 495424
rect 573462 494448 573496 495424
rect 573720 494448 573754 495424
rect 573978 494448 574012 495424
rect 574236 494448 574270 495424
rect 574494 494448 574528 495424
rect 574752 494448 574786 495424
rect 575010 494448 575044 495424
rect 575268 494448 575302 495424
rect 575526 494448 575560 495424
rect 575784 494448 575818 495424
rect 576042 494448 576076 495424
rect 576300 494448 576334 495424
rect 576558 494448 576592 495424
rect 576816 494448 576850 495424
rect 577074 494448 577108 495424
rect 577332 494448 577366 495424
rect 577590 494448 577624 495424
rect 577704 494418 577738 495392
rect 572534 494364 572618 494398
rect 572792 494364 572876 494398
rect 573050 494364 573134 494398
rect 573308 494364 573392 494398
rect 573566 494364 573650 494398
rect 573824 494364 573908 494398
rect 574082 494364 574166 494398
rect 574340 494364 574424 494398
rect 574598 494364 574682 494398
rect 574856 494364 574940 494398
rect 575114 494364 575198 494398
rect 575372 494364 575456 494398
rect 575630 494364 575714 494398
rect 575888 494364 575972 494398
rect 576146 494364 576230 494398
rect 576404 494364 576488 494398
rect 576662 494364 576746 494398
rect 576920 494364 577004 494398
rect 577178 494364 577262 494398
rect 577436 494364 577520 494398
rect 503920 475284 504020 475306
rect 504144 475284 504244 475306
rect 504368 475284 504468 475306
rect 504592 475284 504692 475306
rect 504816 475284 504916 475306
rect 505040 475284 505140 475306
rect 505264 475284 505364 475306
rect 505488 475284 505588 475306
rect 505712 475284 505812 475306
rect 505936 475284 506036 475306
rect 506160 475284 506260 475306
rect 506384 475284 506484 475306
rect 506608 475284 506708 475306
rect 506832 475284 506932 475306
rect 507056 475284 507156 475306
rect 507280 475284 507380 475306
rect 507504 475284 507604 475306
rect 507728 475284 507828 475306
rect 507952 475284 508052 475306
rect 508176 475284 508276 475306
rect 508400 475284 508500 475306
rect 508624 475284 508724 475306
rect 508848 475284 508948 475306
rect 509072 475284 509172 475306
rect 509296 475284 509396 475306
rect 509520 475284 509620 475306
rect 509744 475284 509844 475306
rect 509968 475284 510068 475306
rect 510192 475284 510292 475306
rect 510416 475284 510516 475306
rect 517320 475284 517420 475306
rect 517544 475284 517644 475306
rect 517768 475284 517868 475306
rect 517992 475284 518092 475306
rect 518216 475284 518316 475306
rect 518440 475284 518540 475306
rect 518664 475284 518764 475306
rect 518888 475284 518988 475306
rect 519112 475284 519212 475306
rect 519336 475284 519436 475306
rect 519560 475284 519660 475306
rect 519784 475284 519884 475306
rect 520008 475284 520108 475306
rect 520232 475284 520332 475306
rect 520456 475284 520556 475306
rect 520680 475284 520780 475306
rect 520904 475284 521004 475306
rect 521128 475284 521228 475306
rect 521352 475284 521452 475306
rect 521576 475284 521676 475306
rect 521800 475284 521900 475306
rect 522024 475284 522124 475306
rect 522248 475284 522348 475306
rect 522472 475284 522572 475306
rect 522696 475284 522796 475306
rect 522920 475284 523020 475306
rect 523144 475284 523244 475306
rect 523368 475284 523468 475306
rect 523592 475284 523692 475306
rect 523816 475284 523916 475306
rect 503920 475206 504020 475284
rect 504144 475206 504244 475284
rect 504368 475206 504468 475284
rect 504592 475206 504692 475284
rect 504816 475206 504916 475284
rect 505040 475206 505140 475284
rect 505264 475206 505364 475284
rect 505488 475206 505588 475284
rect 505712 475206 505812 475284
rect 505936 475206 506036 475284
rect 506160 475206 506260 475284
rect 506384 475206 506484 475284
rect 506608 475206 506708 475284
rect 506832 475206 506932 475284
rect 507056 475206 507156 475284
rect 507280 475206 507380 475284
rect 507504 475206 507604 475284
rect 507728 475206 507828 475284
rect 507952 475206 508052 475284
rect 508176 475206 508276 475284
rect 508400 475206 508500 475284
rect 508624 475206 508724 475284
rect 508848 475206 508948 475284
rect 509072 475206 509172 475284
rect 509296 475206 509396 475284
rect 509520 475206 509620 475284
rect 509744 475206 509844 475284
rect 509968 475206 510068 475284
rect 510192 475206 510292 475284
rect 510416 475206 510516 475284
rect 517320 475206 517420 475284
rect 517544 475206 517644 475284
rect 517768 475206 517868 475284
rect 517992 475206 518092 475284
rect 518216 475206 518316 475284
rect 518440 475206 518540 475284
rect 518664 475206 518764 475284
rect 518888 475206 518988 475284
rect 519112 475206 519212 475284
rect 519336 475206 519436 475284
rect 519560 475206 519660 475284
rect 519784 475206 519884 475284
rect 520008 475206 520108 475284
rect 520232 475206 520332 475284
rect 520456 475206 520556 475284
rect 520680 475206 520780 475284
rect 520904 475206 521004 475284
rect 521128 475206 521228 475284
rect 521352 475206 521452 475284
rect 521576 475206 521676 475284
rect 521800 475206 521900 475284
rect 522024 475206 522124 475284
rect 522248 475206 522348 475284
rect 522472 475206 522572 475284
rect 522696 475206 522796 475284
rect 522920 475206 523020 475284
rect 523144 475206 523244 475284
rect 523368 475206 523468 475284
rect 523592 475206 523692 475284
rect 523816 475206 523916 475284
rect 503920 474982 504020 475082
rect 504144 474982 504244 475082
rect 504368 474982 504468 475082
rect 504592 474982 504692 475082
rect 504816 474982 504916 475082
rect 505040 474982 505140 475082
rect 505264 474982 505364 475082
rect 505488 474982 505588 475082
rect 505712 474982 505812 475082
rect 505936 474982 506036 475082
rect 506160 474982 506260 475082
rect 506384 474982 506484 475082
rect 506608 474982 506708 475082
rect 506832 474982 506932 475082
rect 507056 474982 507156 475082
rect 507280 474982 507380 475082
rect 507504 474982 507604 475082
rect 507728 474982 507828 475082
rect 507952 474982 508052 475082
rect 508176 474982 508276 475082
rect 508400 474982 508500 475082
rect 508624 474982 508724 475082
rect 508848 474982 508948 475082
rect 509072 474982 509172 475082
rect 509296 474982 509396 475082
rect 509520 474982 509620 475082
rect 509744 474982 509844 475082
rect 509968 474982 510068 475082
rect 510192 474982 510292 475082
rect 510416 474982 510516 475082
rect 517320 474982 517420 475082
rect 517544 474982 517644 475082
rect 517768 474982 517868 475082
rect 517992 474982 518092 475082
rect 518216 474982 518316 475082
rect 518440 474982 518540 475082
rect 518664 474982 518764 475082
rect 518888 474982 518988 475082
rect 519112 474982 519212 475082
rect 519336 474982 519436 475082
rect 519560 474982 519660 475082
rect 519784 474982 519884 475082
rect 520008 474982 520108 475082
rect 520232 474982 520332 475082
rect 520456 474982 520556 475082
rect 520680 474982 520780 475082
rect 520904 474982 521004 475082
rect 521128 474982 521228 475082
rect 521352 474982 521452 475082
rect 521576 474982 521676 475082
rect 521800 474982 521900 475082
rect 522024 474982 522124 475082
rect 522248 474982 522348 475082
rect 522472 474982 522572 475082
rect 522696 474982 522796 475082
rect 522920 474982 523020 475082
rect 523144 474982 523244 475082
rect 523368 474982 523468 475082
rect 523592 474982 523692 475082
rect 523816 474982 523916 475082
rect 503920 474758 504020 474858
rect 504144 474758 504244 474858
rect 504368 474758 504468 474858
rect 504592 474758 504692 474858
rect 504816 474758 504916 474858
rect 505040 474758 505140 474858
rect 505264 474758 505364 474858
rect 505488 474758 505588 474858
rect 505712 474758 505812 474858
rect 505936 474758 506036 474858
rect 506160 474758 506260 474858
rect 506384 474758 506484 474858
rect 506608 474758 506708 474858
rect 506832 474758 506932 474858
rect 507056 474758 507156 474858
rect 507280 474758 507380 474858
rect 507504 474758 507604 474858
rect 507728 474758 507828 474858
rect 507952 474758 508052 474858
rect 508176 474758 508276 474858
rect 508400 474758 508500 474858
rect 508624 474758 508724 474858
rect 508848 474758 508948 474858
rect 509072 474758 509172 474858
rect 509296 474758 509396 474858
rect 509520 474758 509620 474858
rect 509744 474758 509844 474858
rect 509968 474758 510068 474858
rect 510192 474758 510292 474858
rect 510416 474758 510516 474858
rect 517320 474758 517420 474858
rect 517544 474758 517644 474858
rect 517768 474758 517868 474858
rect 517992 474758 518092 474858
rect 518216 474758 518316 474858
rect 518440 474758 518540 474858
rect 518664 474758 518764 474858
rect 518888 474758 518988 474858
rect 519112 474758 519212 474858
rect 519336 474758 519436 474858
rect 519560 474758 519660 474858
rect 519784 474758 519884 474858
rect 520008 474758 520108 474858
rect 520232 474758 520332 474858
rect 520456 474758 520556 474858
rect 520680 474758 520780 474858
rect 520904 474758 521004 474858
rect 521128 474758 521228 474858
rect 521352 474758 521452 474858
rect 521576 474758 521676 474858
rect 521800 474758 521900 474858
rect 522024 474758 522124 474858
rect 522248 474758 522348 474858
rect 522472 474758 522572 474858
rect 522696 474758 522796 474858
rect 522920 474758 523020 474858
rect 523144 474758 523244 474858
rect 523368 474758 523468 474858
rect 523592 474758 523692 474858
rect 523816 474758 523916 474858
rect 503920 474534 504020 474634
rect 504144 474534 504244 474634
rect 504368 474534 504468 474634
rect 504592 474534 504692 474634
rect 504816 474534 504916 474634
rect 505040 474534 505140 474634
rect 505264 474534 505364 474634
rect 505488 474534 505588 474634
rect 505712 474534 505812 474634
rect 505936 474534 506036 474634
rect 506160 474534 506260 474634
rect 506384 474534 506484 474634
rect 506608 474534 506708 474634
rect 506832 474534 506932 474634
rect 507056 474534 507156 474634
rect 507280 474534 507380 474634
rect 507504 474534 507604 474634
rect 507728 474534 507828 474634
rect 507952 474534 508052 474634
rect 508176 474534 508276 474634
rect 508400 474534 508500 474634
rect 508624 474534 508724 474634
rect 508848 474534 508948 474634
rect 509072 474534 509172 474634
rect 509296 474534 509396 474634
rect 509520 474534 509620 474634
rect 509744 474534 509844 474634
rect 509968 474534 510068 474634
rect 510192 474534 510292 474634
rect 510416 474534 510516 474634
rect 517320 474534 517420 474634
rect 517544 474534 517644 474634
rect 517768 474534 517868 474634
rect 517992 474534 518092 474634
rect 518216 474534 518316 474634
rect 518440 474534 518540 474634
rect 518664 474534 518764 474634
rect 518888 474534 518988 474634
rect 519112 474534 519212 474634
rect 519336 474534 519436 474634
rect 519560 474534 519660 474634
rect 519784 474534 519884 474634
rect 520008 474534 520108 474634
rect 520232 474534 520332 474634
rect 520456 474534 520556 474634
rect 520680 474534 520780 474634
rect 520904 474534 521004 474634
rect 521128 474534 521228 474634
rect 521352 474534 521452 474634
rect 521576 474534 521676 474634
rect 521800 474534 521900 474634
rect 522024 474534 522124 474634
rect 522248 474534 522348 474634
rect 522472 474534 522572 474634
rect 522696 474534 522796 474634
rect 522920 474534 523020 474634
rect 523144 474534 523244 474634
rect 523368 474534 523468 474634
rect 523592 474534 523692 474634
rect 523816 474534 523916 474634
rect 503920 474310 504020 474410
rect 504144 474310 504244 474410
rect 504368 474310 504468 474410
rect 504592 474310 504692 474410
rect 504816 474310 504916 474410
rect 505040 474310 505140 474410
rect 505264 474310 505364 474410
rect 505488 474310 505588 474410
rect 505712 474310 505812 474410
rect 505936 474310 506036 474410
rect 506160 474310 506260 474410
rect 506384 474310 506484 474410
rect 506608 474310 506708 474410
rect 506832 474310 506932 474410
rect 507056 474310 507156 474410
rect 507280 474310 507380 474410
rect 507504 474310 507604 474410
rect 507728 474310 507828 474410
rect 507952 474310 508052 474410
rect 508176 474310 508276 474410
rect 508400 474310 508500 474410
rect 508624 474310 508724 474410
rect 508848 474310 508948 474410
rect 509072 474310 509172 474410
rect 509296 474310 509396 474410
rect 509520 474310 509620 474410
rect 509744 474310 509844 474410
rect 509968 474310 510068 474410
rect 510192 474310 510292 474410
rect 510416 474310 510516 474410
rect 517320 474310 517420 474410
rect 517544 474310 517644 474410
rect 517768 474310 517868 474410
rect 517992 474310 518092 474410
rect 518216 474310 518316 474410
rect 518440 474310 518540 474410
rect 518664 474310 518764 474410
rect 518888 474310 518988 474410
rect 519112 474310 519212 474410
rect 519336 474310 519436 474410
rect 519560 474310 519660 474410
rect 519784 474310 519884 474410
rect 520008 474310 520108 474410
rect 520232 474310 520332 474410
rect 520456 474310 520556 474410
rect 520680 474310 520780 474410
rect 520904 474310 521004 474410
rect 521128 474310 521228 474410
rect 521352 474310 521452 474410
rect 521576 474310 521676 474410
rect 521800 474310 521900 474410
rect 522024 474310 522124 474410
rect 522248 474310 522348 474410
rect 522472 474310 522572 474410
rect 522696 474310 522796 474410
rect 522920 474310 523020 474410
rect 523144 474310 523244 474410
rect 523368 474310 523468 474410
rect 523592 474310 523692 474410
rect 523816 474310 523916 474410
rect 500398 474180 500498 474280
rect 500622 474180 500722 474280
rect 500846 474180 500946 474280
rect 501070 474180 501170 474280
rect 501294 474180 501368 474280
rect 501368 474180 501394 474280
rect 500398 473956 500498 474056
rect 500622 473956 500722 474056
rect 500846 473956 500946 474056
rect 501070 473956 501170 474056
rect 501294 473956 501368 474056
rect 501368 473956 501394 474056
rect 500398 473732 500498 473832
rect 500622 473732 500722 473832
rect 500846 473732 500946 473832
rect 501070 473732 501170 473832
rect 501294 473732 501368 473832
rect 501368 473732 501394 473832
rect 500398 473508 500498 473608
rect 500622 473508 500722 473608
rect 500846 473508 500946 473608
rect 501070 473508 501170 473608
rect 501294 473508 501368 473608
rect 501368 473508 501394 473608
rect 500398 473284 500498 473384
rect 500622 473284 500722 473384
rect 500846 473284 500946 473384
rect 501070 473284 501170 473384
rect 501294 473284 501368 473384
rect 501368 473284 501394 473384
rect 500398 473060 500498 473160
rect 500622 473060 500722 473160
rect 500846 473060 500946 473160
rect 501070 473060 501170 473160
rect 501294 473060 501368 473160
rect 501368 473060 501394 473160
rect 500398 472836 500498 472936
rect 500622 472836 500722 472936
rect 500846 472836 500946 472936
rect 501070 472836 501170 472936
rect 501294 472836 501368 472936
rect 501368 472836 501394 472936
rect 506570 472730 506946 472764
rect 500398 472612 500498 472712
rect 500622 472612 500722 472712
rect 500846 472612 500946 472712
rect 501070 472612 501170 472712
rect 501294 472612 501368 472712
rect 501368 472612 501394 472712
rect 500398 472388 500498 472488
rect 500622 472388 500722 472488
rect 500846 472388 500946 472488
rect 501070 472388 501170 472488
rect 501294 472388 501368 472488
rect 501368 472388 501394 472488
rect 506996 472426 507030 472610
rect 525680 472468 526478 472484
rect 506570 472272 506946 472306
rect 500398 472164 500498 472264
rect 500622 472164 500722 472264
rect 500846 472164 500946 472264
rect 501070 472164 501170 472264
rect 501294 472164 501368 472264
rect 501368 472164 501394 472264
rect 500398 471940 500498 472040
rect 500622 471940 500722 472040
rect 500846 471940 500946 472040
rect 501070 471940 501170 472040
rect 501294 471940 501368 472040
rect 501368 471940 501394 472040
rect 506996 471968 507030 472152
rect 500398 471716 500498 471816
rect 500622 471716 500722 471816
rect 500846 471716 500946 471816
rect 501070 471716 501170 471816
rect 501294 471716 501368 471816
rect 501368 471716 501394 471816
rect 506570 471814 506946 471848
rect 500398 471492 500498 471592
rect 500622 471492 500722 471592
rect 500846 471492 500946 471592
rect 501070 471492 501170 471592
rect 501294 471492 501368 471592
rect 501368 471492 501394 471592
rect 506996 471510 507030 471694
rect 500398 471268 500498 471368
rect 500622 471268 500722 471368
rect 500846 471268 500946 471368
rect 501070 471268 501170 471368
rect 501294 471268 501368 471368
rect 501368 471268 501394 471368
rect 506570 471356 506946 471390
rect 500398 471044 500498 471144
rect 500622 471044 500722 471144
rect 500846 471044 500946 471144
rect 501070 471044 501170 471144
rect 501294 471044 501368 471144
rect 501368 471044 501394 471144
rect 506996 471052 507030 471236
rect 500398 470820 500498 470920
rect 500622 470820 500722 470920
rect 500846 470820 500946 470920
rect 501070 470820 501170 470920
rect 501294 470820 501368 470920
rect 501368 470820 501394 470920
rect 506570 470898 506946 470932
rect 507094 471806 507146 471858
rect 507094 470890 507146 470942
rect 500398 470596 500498 470696
rect 500622 470596 500722 470696
rect 500846 470596 500946 470696
rect 501070 470596 501170 470696
rect 501294 470596 501368 470696
rect 501368 470596 501394 470696
rect 506996 470594 507030 470778
rect 500398 470372 500498 470472
rect 500622 470372 500722 470472
rect 500846 470372 500946 470472
rect 501070 470372 501170 470472
rect 501294 470372 501368 470472
rect 501368 470372 501394 470472
rect 506570 470440 506946 470474
rect 500398 470148 500498 470248
rect 500622 470148 500722 470248
rect 500846 470148 500946 470248
rect 501070 470148 501170 470248
rect 501294 470148 501368 470248
rect 501368 470148 501394 470248
rect 503226 470102 505568 470202
rect 506996 470136 507030 470320
rect 500398 469924 500498 470024
rect 500622 469924 500722 470024
rect 500846 469924 500946 470024
rect 501070 469924 501170 470024
rect 501294 469924 501368 470024
rect 501368 469924 501394 470024
rect 506570 469982 506946 470016
rect 500398 469700 500498 469800
rect 500622 469700 500722 469800
rect 500846 469700 500946 469800
rect 501070 469700 501170 469800
rect 501294 469700 501368 469800
rect 501368 469700 501394 469800
rect 500398 469476 500498 469576
rect 500622 469476 500722 469576
rect 500846 469476 500946 469576
rect 501070 469476 501170 469576
rect 501294 469476 501368 469576
rect 501368 469476 501394 469576
rect 503100 469526 505656 469560
rect 500398 469252 500498 469352
rect 500622 469252 500722 469352
rect 500846 469252 500946 469352
rect 501070 469252 501170 469352
rect 501294 469252 501368 469352
rect 501368 469252 501394 469352
rect 505715 469222 505749 469406
rect 500398 469028 500498 469128
rect 500622 469028 500722 469128
rect 500846 469028 500946 469128
rect 501070 469028 501170 469128
rect 501294 469028 501368 469128
rect 501368 469028 501394 469128
rect 503100 469068 505656 469102
rect 503100 468954 505656 468988
rect 500398 468804 500498 468904
rect 500622 468804 500722 468904
rect 500846 468804 500946 468904
rect 501070 468804 501170 468904
rect 501294 468804 501368 468904
rect 501368 468804 501394 468904
rect 500398 468580 500498 468680
rect 500622 468580 500722 468680
rect 500846 468580 500946 468680
rect 501070 468580 501170 468680
rect 501294 468580 501368 468680
rect 501368 468580 501394 468680
rect 505715 468650 505749 468834
rect 503100 468496 505656 468530
rect 500398 468356 500498 468456
rect 500622 468356 500722 468456
rect 500846 468356 500946 468456
rect 501070 468356 501170 468456
rect 501294 468356 501368 468456
rect 501368 468356 501394 468456
rect 503100 468382 505656 468416
rect 506470 468286 508068 468386
rect 500398 468132 500498 468232
rect 500622 468132 500722 468232
rect 500846 468132 500946 468232
rect 501070 468132 501170 468232
rect 501294 468132 501368 468232
rect 501368 468132 501394 468232
rect 505715 468078 505749 468262
rect 509940 468166 510124 468200
rect 500398 467908 500498 468008
rect 500622 467908 500722 468008
rect 500846 467908 500946 468008
rect 501070 467908 501170 468008
rect 501294 467908 501368 468008
rect 501368 467908 501394 468008
rect 503100 467924 505656 467958
rect 503100 467810 505656 467844
rect 506292 467800 508068 467834
rect 500398 467684 500498 467784
rect 500622 467684 500722 467784
rect 500846 467684 500946 467784
rect 501070 467684 501170 467784
rect 501294 467684 501368 467784
rect 501368 467684 501394 467784
rect 505715 467506 505749 467690
rect 508118 467496 508152 467680
rect 503100 467352 505656 467386
rect 506292 467342 508068 467376
rect 503100 467238 505656 467272
rect 506292 467228 508068 467262
rect 505715 466934 505749 467118
rect 508118 466924 508152 467108
rect 503100 466780 505656 466814
rect 506292 466770 508068 466804
rect 503100 466666 505656 466700
rect 506292 466656 508068 466690
rect 502622 464278 502722 466620
rect 505715 466362 505749 466546
rect 508118 466352 508152 466536
rect 503100 466208 505656 466242
rect 506292 466198 508068 466232
rect 503100 466094 505656 466128
rect 506292 466084 508068 466118
rect 505715 465790 505749 465974
rect 508118 465780 508152 465964
rect 503100 465636 505656 465670
rect 506292 465626 508068 465660
rect 503100 465522 505656 465556
rect 506292 465512 508068 465546
rect 505715 465218 505749 465402
rect 508118 465208 508152 465392
rect 503100 465064 505656 465098
rect 506292 465054 508068 465088
rect 503100 464950 505656 464984
rect 506292 464940 508068 464974
rect 505715 464646 505749 464830
rect 508118 464636 508152 464820
rect 503100 464492 505656 464526
rect 506292 464482 508068 464516
rect 503100 464378 505656 464412
rect 506292 464368 508068 464402
rect 505715 464074 505749 464258
rect 508118 464064 508152 464248
rect 503100 463920 505656 463954
rect 506292 463910 508068 463944
rect 500398 463710 500498 463810
rect 500622 463710 500722 463810
rect 500846 463710 500946 463810
rect 501070 463710 501170 463810
rect 501294 463710 501368 463810
rect 501368 463710 501394 463810
rect 503100 463806 505656 463840
rect 506292 463796 508068 463830
rect 500398 463486 500498 463586
rect 500622 463486 500722 463586
rect 500846 463486 500946 463586
rect 501070 463486 501170 463586
rect 501294 463486 501368 463586
rect 501368 463486 501394 463586
rect 505715 463502 505749 463686
rect 508118 463492 508152 463676
rect 500398 463262 500498 463362
rect 500622 463262 500722 463362
rect 500846 463262 500946 463362
rect 501070 463262 501170 463362
rect 501294 463262 501368 463362
rect 501368 463262 501394 463362
rect 503100 463348 505656 463382
rect 506292 463338 508068 463372
rect 503100 463234 505656 463268
rect 500398 463038 500498 463138
rect 500622 463038 500722 463138
rect 500846 463038 500946 463138
rect 501070 463038 501170 463138
rect 501294 463038 501368 463138
rect 501368 463038 501394 463138
rect 505715 462930 505749 463114
rect 500398 462814 500498 462914
rect 500622 462814 500722 462914
rect 500846 462814 500946 462914
rect 501070 462814 501170 462914
rect 501294 462814 501368 462914
rect 501368 462814 501394 462914
rect 503100 462776 505656 462810
rect 506470 462786 508068 462886
rect 509786 462740 509820 468116
rect 510244 462740 510278 468116
rect 500398 462590 500498 462690
rect 500622 462590 500722 462690
rect 500846 462590 500946 462690
rect 501070 462590 501170 462690
rect 501294 462590 501368 462690
rect 501368 462590 501394 462690
rect 503100 462662 505656 462696
rect 500398 462366 500498 462466
rect 500622 462366 500722 462466
rect 500846 462366 500946 462466
rect 501070 462366 501170 462466
rect 501294 462366 501368 462466
rect 501368 462366 501394 462466
rect 505715 462358 505749 462542
rect 510470 468834 510814 468840
rect 510470 462382 510476 468834
rect 510476 462382 510808 468834
rect 510808 462382 510814 468834
rect 510470 462376 510814 462382
rect 500398 462142 500498 462242
rect 500622 462142 500722 462242
rect 500846 462142 500946 462242
rect 501070 462142 501170 462242
rect 501294 462142 501368 462242
rect 501368 462142 501394 462242
rect 503100 462204 505656 462238
rect 503100 462090 505656 462124
rect 500398 461918 500498 462018
rect 500622 461918 500722 462018
rect 500846 461918 500946 462018
rect 501070 461918 501170 462018
rect 501294 461918 501368 462018
rect 501368 461918 501394 462018
rect 500398 461694 500498 461794
rect 500622 461694 500722 461794
rect 500846 461694 500946 461794
rect 501070 461694 501170 461794
rect 501294 461694 501368 461794
rect 501368 461694 501394 461794
rect 505715 461786 505749 461970
rect 503100 461632 505656 461666
rect 500398 461470 500498 461570
rect 500622 461470 500722 461570
rect 500846 461470 500946 461570
rect 501070 461470 501170 461570
rect 501294 461470 501368 461570
rect 501368 461470 501394 461570
rect 500398 461246 500498 461346
rect 500622 461246 500722 461346
rect 500846 461246 500946 461346
rect 501070 461246 501170 461346
rect 501294 461246 501368 461346
rect 501368 461246 501394 461346
rect 525680 461284 525696 472468
rect 525696 461284 526462 472468
rect 526462 461284 526478 472468
rect 525680 461268 526478 461284
rect 500398 461022 500498 461122
rect 500622 461022 500722 461122
rect 500846 461022 500946 461122
rect 501070 461022 501170 461122
rect 501294 461022 501368 461122
rect 501368 461022 501394 461122
rect 503226 460974 505568 461074
rect 500398 460798 500498 460898
rect 500622 460798 500722 460898
rect 500846 460798 500946 460898
rect 501070 460798 501170 460898
rect 501294 460798 501368 460898
rect 501368 460798 501394 460898
rect 500398 460574 500498 460674
rect 500622 460574 500722 460674
rect 500846 460574 500946 460674
rect 501070 460574 501170 460674
rect 501294 460574 501368 460674
rect 501368 460574 501394 460674
rect 500398 460350 500498 460450
rect 500622 460350 500722 460450
rect 500846 460350 500946 460450
rect 501070 460350 501170 460450
rect 501294 460350 501368 460450
rect 501368 460350 501394 460450
rect 500398 460126 500498 460226
rect 500622 460126 500722 460226
rect 500846 460126 500946 460226
rect 501070 460126 501170 460226
rect 501294 460126 501368 460226
rect 501368 460126 501394 460226
rect 500398 459902 500498 460002
rect 500622 459902 500722 460002
rect 500846 459902 500946 460002
rect 501070 459902 501170 460002
rect 501294 459902 501368 460002
rect 501368 459902 501394 460002
rect 502528 459952 502628 460352
rect 500398 459678 500498 459778
rect 500622 459678 500722 459778
rect 500846 459678 500946 459778
rect 501070 459678 501170 459778
rect 501294 459678 501368 459778
rect 501368 459678 501394 459778
rect 503138 459718 510854 459752
rect 500398 459454 500498 459554
rect 500622 459454 500722 459554
rect 500846 459454 500946 459554
rect 501070 459454 501170 459554
rect 501294 459454 501368 459554
rect 501368 459454 501394 459554
rect 503045 459414 503079 459598
rect 500398 459230 500498 459330
rect 500622 459230 500722 459330
rect 500846 459230 500946 459330
rect 501070 459230 501170 459330
rect 501294 459230 501368 459330
rect 501368 459230 501394 459330
rect 517864 459330 518261 459868
rect 521619 459330 522016 459868
rect 503138 459260 510854 459294
rect 500398 459006 500498 459106
rect 500622 459006 500722 459106
rect 500846 459006 500946 459106
rect 501070 459006 501170 459106
rect 501294 459006 501368 459106
rect 501368 459006 501394 459106
rect 503045 458956 503079 459140
rect 500398 458782 500498 458882
rect 500622 458782 500722 458882
rect 500846 458782 500946 458882
rect 501070 458782 501170 458882
rect 501294 458782 501368 458882
rect 501368 458782 501394 458882
rect 503138 458802 510854 458836
rect 500398 458558 500498 458658
rect 500622 458558 500722 458658
rect 500846 458558 500946 458658
rect 501070 458558 501170 458658
rect 501294 458558 501368 458658
rect 501368 458558 501394 458658
rect 503045 458498 503079 458682
rect 500398 458334 500498 458434
rect 500622 458334 500722 458434
rect 500846 458334 500946 458434
rect 501070 458334 501170 458434
rect 501294 458334 501368 458434
rect 501368 458334 501394 458434
rect 503138 458344 510854 458378
rect 500398 458110 500498 458210
rect 500622 458110 500722 458210
rect 500846 458110 500946 458210
rect 501070 458110 501170 458210
rect 501294 458110 501368 458210
rect 501368 458110 501394 458210
rect 503045 458040 503079 458224
rect 500398 457886 500498 457986
rect 500622 457886 500722 457986
rect 500846 457886 500946 457986
rect 501070 457886 501170 457986
rect 501294 457886 501368 457986
rect 501368 457886 501394 457986
rect 503138 457886 510854 457920
rect 500398 457662 500498 457762
rect 500622 457662 500722 457762
rect 500846 457662 500946 457762
rect 501070 457662 501170 457762
rect 501294 457662 501368 457762
rect 501368 457662 501394 457762
rect 503045 457582 503079 457766
rect 500398 457438 500498 457538
rect 500622 457438 500722 457538
rect 500846 457438 500946 457538
rect 501070 457438 501170 457538
rect 501294 457438 501368 457538
rect 501368 457438 501394 457538
rect 517864 458512 518261 459050
rect 521619 458512 522016 459050
rect 517864 457694 518261 458232
rect 521619 457694 522016 458232
rect 503138 457428 510854 457462
rect 500398 457214 500498 457314
rect 500622 457214 500722 457314
rect 500846 457214 500946 457314
rect 501070 457214 501170 457314
rect 501294 457214 501368 457314
rect 501368 457214 501394 457314
rect 503045 457124 503079 457308
rect 503138 456970 510854 457004
rect 517594 456918 518660 457412
rect 503045 456666 503079 456850
rect 503138 456512 510854 456546
rect 503045 456208 503079 456392
rect 503138 456054 510854 456088
rect 518274 456058 518671 456596
rect 523005 456058 523402 456596
rect 503045 455750 503079 455934
rect 503138 455596 510854 455630
rect 503045 455292 503079 455476
rect 518274 455240 518671 455778
rect 523005 455240 523402 455778
rect 503138 455138 510854 455172
rect 503045 454834 503079 455018
rect 503138 454680 510854 454714
rect 502528 454042 502628 454442
rect 518274 454422 518671 454960
rect 523005 454422 523402 454960
rect 503138 453760 510854 453794
rect 503045 453456 503079 453640
rect 518274 453604 518671 454142
rect 503138 453302 510854 453336
rect 503045 452998 503079 453182
rect 503138 452844 510854 452878
rect 503045 452540 503079 452724
rect 523005 453604 523402 454142
rect 503138 452386 510854 452420
rect 503045 452082 503079 452266
rect 503138 451928 510854 451962
rect 517606 451948 518658 452460
rect 503045 451624 503079 451808
rect 503138 451470 510854 451504
rect 503045 451166 503079 451350
rect 516208 451150 516605 451688
rect 522943 451150 523340 451688
rect 503138 451012 510854 451046
rect 503045 450708 503079 450892
rect 503138 450554 510854 450588
rect 503045 450250 503079 450434
rect 516207 450332 516605 450870
rect 522943 450332 523340 450870
rect 503138 450096 510854 450130
rect 503045 449792 503079 449976
rect 503138 449638 510854 449672
rect 503045 449334 503079 449518
rect 516208 449514 516605 450052
rect 522943 449514 523340 450052
rect 503138 449180 510854 449214
rect 502528 448542 502628 448942
rect 516208 448696 516605 449234
rect 522943 448696 523340 449234
rect 503138 448260 510854 448294
rect 503045 447956 503079 448140
rect 516207 447878 516605 448416
rect 522943 447878 523340 448416
rect 503138 447802 510854 447836
rect 503045 447498 503079 447682
rect 503138 447344 510854 447378
rect 503045 447040 503079 447224
rect 516208 447060 516605 447598
rect 522943 447060 523340 447598
rect 503138 446886 510854 446920
rect 503045 446582 503079 446766
rect 503138 446428 510854 446462
rect 503045 446124 503079 446308
rect 516208 446242 516605 446780
rect 522943 446242 523340 446780
rect 503138 445970 510854 446004
rect 503045 445666 503079 445850
rect 503138 445512 510854 445546
rect 516207 445424 516605 445962
rect 522943 445424 523340 445962
rect 503045 445208 503079 445392
rect 503138 445054 510854 445088
rect 503045 444750 503079 444934
rect 503138 444596 510854 444630
rect 516208 444606 516605 445144
rect 522943 444606 523340 445144
rect 503045 444292 503079 444476
rect 503138 444138 510854 444172
rect 503045 443834 503079 444018
rect 516208 443788 516605 444326
rect 522943 443788 523340 444326
rect 503138 443680 510854 443714
rect 503045 443376 503079 443560
rect 503138 443222 510854 443256
rect 502526 442586 502626 442986
rect 516208 442970 516605 443508
rect 522943 442970 523340 443508
rect 516207 442152 516605 442690
rect 522943 442152 523340 442690
rect 516208 441334 516605 441872
rect 522943 441334 523340 441872
rect 516208 440516 516605 441054
rect 522943 440516 523340 441054
rect 516208 439698 516605 440236
rect 522943 439698 523340 440236
rect 516208 438880 516605 439418
rect 522943 438880 523340 439418
rect 500418 437440 500518 437540
rect 500642 437440 500742 437540
rect 500866 437440 500966 437540
rect 501090 437440 501190 437540
rect 501314 437440 501368 437540
rect 501368 437440 501414 437540
rect 503740 438090 503762 438112
rect 503762 438090 503774 438112
rect 503840 438090 503852 438112
rect 503852 438090 503874 438112
rect 503940 438090 503942 438112
rect 503942 438090 503974 438112
rect 503740 438078 503774 438090
rect 503840 438078 503874 438090
rect 503940 438078 503974 438090
rect 504040 438078 504074 438112
rect 504140 438078 504174 438112
rect 504240 438090 504268 438112
rect 504268 438090 504274 438112
rect 504240 438078 504274 438090
rect 503740 438000 503762 438012
rect 503762 438000 503774 438012
rect 503840 438000 503852 438012
rect 503852 438000 503874 438012
rect 503940 438000 503942 438012
rect 503942 438000 503974 438012
rect 503740 437978 503774 438000
rect 503840 437978 503874 438000
rect 503940 437978 503974 438000
rect 504040 437978 504074 438012
rect 504140 437978 504174 438012
rect 504240 438000 504268 438012
rect 504268 438000 504274 438012
rect 504240 437978 504274 438000
rect 503740 437910 503762 437912
rect 503762 437910 503774 437912
rect 503840 437910 503852 437912
rect 503852 437910 503874 437912
rect 503940 437910 503942 437912
rect 503942 437910 503974 437912
rect 503740 437878 503774 437910
rect 503840 437878 503874 437910
rect 503940 437878 503974 437910
rect 504040 437878 504074 437912
rect 504140 437878 504174 437912
rect 504240 437910 504268 437912
rect 504268 437910 504274 437912
rect 504240 437878 504274 437910
rect 503740 437778 503774 437812
rect 503840 437778 503874 437812
rect 503940 437778 503974 437812
rect 504040 437778 504074 437812
rect 504140 437778 504174 437812
rect 504240 437778 504274 437812
rect 503740 437678 503774 437712
rect 503840 437678 503874 437712
rect 503940 437678 503974 437712
rect 504040 437678 504074 437712
rect 504140 437678 504174 437712
rect 504240 437678 504274 437712
rect 503740 437584 503774 437612
rect 503840 437584 503874 437612
rect 503940 437584 503974 437612
rect 503740 437578 503762 437584
rect 503762 437578 503774 437584
rect 503840 437578 503852 437584
rect 503852 437578 503874 437584
rect 503940 437578 503942 437584
rect 503942 437578 503974 437584
rect 504040 437578 504074 437612
rect 504140 437578 504174 437612
rect 504240 437584 504274 437612
rect 504240 437578 504268 437584
rect 504268 437578 504274 437584
rect 505028 438090 505050 438112
rect 505050 438090 505062 438112
rect 505128 438090 505140 438112
rect 505140 438090 505162 438112
rect 505228 438090 505230 438112
rect 505230 438090 505262 438112
rect 505028 438078 505062 438090
rect 505128 438078 505162 438090
rect 505228 438078 505262 438090
rect 505328 438078 505362 438112
rect 505428 438078 505462 438112
rect 505528 438090 505556 438112
rect 505556 438090 505562 438112
rect 505528 438078 505562 438090
rect 505028 438000 505050 438012
rect 505050 438000 505062 438012
rect 505128 438000 505140 438012
rect 505140 438000 505162 438012
rect 505228 438000 505230 438012
rect 505230 438000 505262 438012
rect 505028 437978 505062 438000
rect 505128 437978 505162 438000
rect 505228 437978 505262 438000
rect 505328 437978 505362 438012
rect 505428 437978 505462 438012
rect 505528 438000 505556 438012
rect 505556 438000 505562 438012
rect 505528 437978 505562 438000
rect 505028 437910 505050 437912
rect 505050 437910 505062 437912
rect 505128 437910 505140 437912
rect 505140 437910 505162 437912
rect 505228 437910 505230 437912
rect 505230 437910 505262 437912
rect 505028 437878 505062 437910
rect 505128 437878 505162 437910
rect 505228 437878 505262 437910
rect 505328 437878 505362 437912
rect 505428 437878 505462 437912
rect 505528 437910 505556 437912
rect 505556 437910 505562 437912
rect 505528 437878 505562 437910
rect 505028 437778 505062 437812
rect 505128 437778 505162 437812
rect 505228 437778 505262 437812
rect 505328 437778 505362 437812
rect 505428 437778 505462 437812
rect 505528 437778 505562 437812
rect 505028 437678 505062 437712
rect 505128 437678 505162 437712
rect 505228 437678 505262 437712
rect 505328 437678 505362 437712
rect 505428 437678 505462 437712
rect 505528 437678 505562 437712
rect 505028 437584 505062 437612
rect 505128 437584 505162 437612
rect 505228 437584 505262 437612
rect 505028 437578 505050 437584
rect 505050 437578 505062 437584
rect 505128 437578 505140 437584
rect 505140 437578 505162 437584
rect 505228 437578 505230 437584
rect 505230 437578 505262 437584
rect 505328 437578 505362 437612
rect 505428 437578 505462 437612
rect 505528 437584 505562 437612
rect 505528 437578 505556 437584
rect 505556 437578 505562 437584
rect 506316 438090 506338 438112
rect 506338 438090 506350 438112
rect 506416 438090 506428 438112
rect 506428 438090 506450 438112
rect 506516 438090 506518 438112
rect 506518 438090 506550 438112
rect 506316 438078 506350 438090
rect 506416 438078 506450 438090
rect 506516 438078 506550 438090
rect 506616 438078 506650 438112
rect 506716 438078 506750 438112
rect 506816 438090 506844 438112
rect 506844 438090 506850 438112
rect 506816 438078 506850 438090
rect 506316 438000 506338 438012
rect 506338 438000 506350 438012
rect 506416 438000 506428 438012
rect 506428 438000 506450 438012
rect 506516 438000 506518 438012
rect 506518 438000 506550 438012
rect 506316 437978 506350 438000
rect 506416 437978 506450 438000
rect 506516 437978 506550 438000
rect 506616 437978 506650 438012
rect 506716 437978 506750 438012
rect 506816 438000 506844 438012
rect 506844 438000 506850 438012
rect 506816 437978 506850 438000
rect 506316 437910 506338 437912
rect 506338 437910 506350 437912
rect 506416 437910 506428 437912
rect 506428 437910 506450 437912
rect 506516 437910 506518 437912
rect 506518 437910 506550 437912
rect 506316 437878 506350 437910
rect 506416 437878 506450 437910
rect 506516 437878 506550 437910
rect 506616 437878 506650 437912
rect 506716 437878 506750 437912
rect 506816 437910 506844 437912
rect 506844 437910 506850 437912
rect 506816 437878 506850 437910
rect 506316 437778 506350 437812
rect 506416 437778 506450 437812
rect 506516 437778 506550 437812
rect 506616 437778 506650 437812
rect 506716 437778 506750 437812
rect 506816 437778 506850 437812
rect 506316 437678 506350 437712
rect 506416 437678 506450 437712
rect 506516 437678 506550 437712
rect 506616 437678 506650 437712
rect 506716 437678 506750 437712
rect 506816 437678 506850 437712
rect 506316 437584 506350 437612
rect 506416 437584 506450 437612
rect 506516 437584 506550 437612
rect 506316 437578 506338 437584
rect 506338 437578 506350 437584
rect 506416 437578 506428 437584
rect 506428 437578 506450 437584
rect 506516 437578 506518 437584
rect 506518 437578 506550 437584
rect 506616 437578 506650 437612
rect 506716 437578 506750 437612
rect 506816 437584 506850 437612
rect 506816 437578 506844 437584
rect 506844 437578 506850 437584
rect 507604 438090 507626 438112
rect 507626 438090 507638 438112
rect 507704 438090 507716 438112
rect 507716 438090 507738 438112
rect 507804 438090 507806 438112
rect 507806 438090 507838 438112
rect 507604 438078 507638 438090
rect 507704 438078 507738 438090
rect 507804 438078 507838 438090
rect 507904 438078 507938 438112
rect 508004 438078 508038 438112
rect 508104 438090 508132 438112
rect 508132 438090 508138 438112
rect 508104 438078 508138 438090
rect 507604 438000 507626 438012
rect 507626 438000 507638 438012
rect 507704 438000 507716 438012
rect 507716 438000 507738 438012
rect 507804 438000 507806 438012
rect 507806 438000 507838 438012
rect 507604 437978 507638 438000
rect 507704 437978 507738 438000
rect 507804 437978 507838 438000
rect 507904 437978 507938 438012
rect 508004 437978 508038 438012
rect 508104 438000 508132 438012
rect 508132 438000 508138 438012
rect 508104 437978 508138 438000
rect 507604 437910 507626 437912
rect 507626 437910 507638 437912
rect 507704 437910 507716 437912
rect 507716 437910 507738 437912
rect 507804 437910 507806 437912
rect 507806 437910 507838 437912
rect 507604 437878 507638 437910
rect 507704 437878 507738 437910
rect 507804 437878 507838 437910
rect 507904 437878 507938 437912
rect 508004 437878 508038 437912
rect 508104 437910 508132 437912
rect 508132 437910 508138 437912
rect 508104 437878 508138 437910
rect 507604 437778 507638 437812
rect 507704 437778 507738 437812
rect 507804 437778 507838 437812
rect 507904 437778 507938 437812
rect 508004 437778 508038 437812
rect 508104 437778 508138 437812
rect 507604 437678 507638 437712
rect 507704 437678 507738 437712
rect 507804 437678 507838 437712
rect 507904 437678 507938 437712
rect 508004 437678 508038 437712
rect 508104 437678 508138 437712
rect 507604 437584 507638 437612
rect 507704 437584 507738 437612
rect 507804 437584 507838 437612
rect 507604 437578 507626 437584
rect 507626 437578 507638 437584
rect 507704 437578 507716 437584
rect 507716 437578 507738 437584
rect 507804 437578 507806 437584
rect 507806 437578 507838 437584
rect 507904 437578 507938 437612
rect 508004 437578 508038 437612
rect 508104 437584 508138 437612
rect 508104 437578 508132 437584
rect 508132 437578 508138 437584
rect 508892 438090 508914 438112
rect 508914 438090 508926 438112
rect 508992 438090 509004 438112
rect 509004 438090 509026 438112
rect 509092 438090 509094 438112
rect 509094 438090 509126 438112
rect 508892 438078 508926 438090
rect 508992 438078 509026 438090
rect 509092 438078 509126 438090
rect 509192 438078 509226 438112
rect 509292 438078 509326 438112
rect 509392 438090 509420 438112
rect 509420 438090 509426 438112
rect 509392 438078 509426 438090
rect 508892 438000 508914 438012
rect 508914 438000 508926 438012
rect 508992 438000 509004 438012
rect 509004 438000 509026 438012
rect 509092 438000 509094 438012
rect 509094 438000 509126 438012
rect 508892 437978 508926 438000
rect 508992 437978 509026 438000
rect 509092 437978 509126 438000
rect 509192 437978 509226 438012
rect 509292 437978 509326 438012
rect 509392 438000 509420 438012
rect 509420 438000 509426 438012
rect 509392 437978 509426 438000
rect 508892 437910 508914 437912
rect 508914 437910 508926 437912
rect 508992 437910 509004 437912
rect 509004 437910 509026 437912
rect 509092 437910 509094 437912
rect 509094 437910 509126 437912
rect 508892 437878 508926 437910
rect 508992 437878 509026 437910
rect 509092 437878 509126 437910
rect 509192 437878 509226 437912
rect 509292 437878 509326 437912
rect 509392 437910 509420 437912
rect 509420 437910 509426 437912
rect 509392 437878 509426 437910
rect 508892 437778 508926 437812
rect 508992 437778 509026 437812
rect 509092 437778 509126 437812
rect 509192 437778 509226 437812
rect 509292 437778 509326 437812
rect 509392 437778 509426 437812
rect 508892 437678 508926 437712
rect 508992 437678 509026 437712
rect 509092 437678 509126 437712
rect 509192 437678 509226 437712
rect 509292 437678 509326 437712
rect 509392 437678 509426 437712
rect 508892 437584 508926 437612
rect 508992 437584 509026 437612
rect 509092 437584 509126 437612
rect 508892 437578 508914 437584
rect 508914 437578 508926 437584
rect 508992 437578 509004 437584
rect 509004 437578 509026 437584
rect 509092 437578 509094 437584
rect 509094 437578 509126 437584
rect 509192 437578 509226 437612
rect 509292 437578 509326 437612
rect 509392 437584 509426 437612
rect 509392 437578 509420 437584
rect 509420 437578 509426 437584
rect 510180 438090 510202 438112
rect 510202 438090 510214 438112
rect 510280 438090 510292 438112
rect 510292 438090 510314 438112
rect 510380 438090 510382 438112
rect 510382 438090 510414 438112
rect 510180 438078 510214 438090
rect 510280 438078 510314 438090
rect 510380 438078 510414 438090
rect 510480 438078 510514 438112
rect 510580 438078 510614 438112
rect 510680 438090 510708 438112
rect 510708 438090 510714 438112
rect 510680 438078 510714 438090
rect 510180 438000 510202 438012
rect 510202 438000 510214 438012
rect 510280 438000 510292 438012
rect 510292 438000 510314 438012
rect 510380 438000 510382 438012
rect 510382 438000 510414 438012
rect 510180 437978 510214 438000
rect 510280 437978 510314 438000
rect 510380 437978 510414 438000
rect 510480 437978 510514 438012
rect 510580 437978 510614 438012
rect 510680 438000 510708 438012
rect 510708 438000 510714 438012
rect 510680 437978 510714 438000
rect 510180 437910 510202 437912
rect 510202 437910 510214 437912
rect 510280 437910 510292 437912
rect 510292 437910 510314 437912
rect 510380 437910 510382 437912
rect 510382 437910 510414 437912
rect 510180 437878 510214 437910
rect 510280 437878 510314 437910
rect 510380 437878 510414 437910
rect 510480 437878 510514 437912
rect 510580 437878 510614 437912
rect 510680 437910 510708 437912
rect 510708 437910 510714 437912
rect 510680 437878 510714 437910
rect 510180 437778 510214 437812
rect 510280 437778 510314 437812
rect 510380 437778 510414 437812
rect 510480 437778 510514 437812
rect 510580 437778 510614 437812
rect 510680 437778 510714 437812
rect 510180 437678 510214 437712
rect 510280 437678 510314 437712
rect 510380 437678 510414 437712
rect 510480 437678 510514 437712
rect 510580 437678 510614 437712
rect 510680 437678 510714 437712
rect 510180 437584 510214 437612
rect 510280 437584 510314 437612
rect 510380 437584 510414 437612
rect 510180 437578 510202 437584
rect 510202 437578 510214 437584
rect 510280 437578 510292 437584
rect 510292 437578 510314 437584
rect 510380 437578 510382 437584
rect 510382 437578 510414 437584
rect 510480 437578 510514 437612
rect 510580 437578 510614 437612
rect 510680 437584 510714 437612
rect 510680 437578 510708 437584
rect 510708 437578 510714 437584
rect 511468 438090 511490 438112
rect 511490 438090 511502 438112
rect 511568 438090 511580 438112
rect 511580 438090 511602 438112
rect 511668 438090 511670 438112
rect 511670 438090 511702 438112
rect 511468 438078 511502 438090
rect 511568 438078 511602 438090
rect 511668 438078 511702 438090
rect 511768 438078 511802 438112
rect 511868 438078 511902 438112
rect 511968 438090 511996 438112
rect 511996 438090 512002 438112
rect 511968 438078 512002 438090
rect 511468 438000 511490 438012
rect 511490 438000 511502 438012
rect 511568 438000 511580 438012
rect 511580 438000 511602 438012
rect 511668 438000 511670 438012
rect 511670 438000 511702 438012
rect 511468 437978 511502 438000
rect 511568 437978 511602 438000
rect 511668 437978 511702 438000
rect 511768 437978 511802 438012
rect 511868 437978 511902 438012
rect 511968 438000 511996 438012
rect 511996 438000 512002 438012
rect 511968 437978 512002 438000
rect 511468 437910 511490 437912
rect 511490 437910 511502 437912
rect 511568 437910 511580 437912
rect 511580 437910 511602 437912
rect 511668 437910 511670 437912
rect 511670 437910 511702 437912
rect 511468 437878 511502 437910
rect 511568 437878 511602 437910
rect 511668 437878 511702 437910
rect 511768 437878 511802 437912
rect 511868 437878 511902 437912
rect 511968 437910 511996 437912
rect 511996 437910 512002 437912
rect 511968 437878 512002 437910
rect 511468 437778 511502 437812
rect 511568 437778 511602 437812
rect 511668 437778 511702 437812
rect 511768 437778 511802 437812
rect 511868 437778 511902 437812
rect 511968 437778 512002 437812
rect 511468 437678 511502 437712
rect 511568 437678 511602 437712
rect 511668 437678 511702 437712
rect 511768 437678 511802 437712
rect 511868 437678 511902 437712
rect 511968 437678 512002 437712
rect 511468 437584 511502 437612
rect 511568 437584 511602 437612
rect 511668 437584 511702 437612
rect 511468 437578 511490 437584
rect 511490 437578 511502 437584
rect 511568 437578 511580 437584
rect 511580 437578 511602 437584
rect 511668 437578 511670 437584
rect 511670 437578 511702 437584
rect 511768 437578 511802 437612
rect 511868 437578 511902 437612
rect 511968 437584 512002 437612
rect 511968 437578 511996 437584
rect 511996 437578 512002 437584
rect 512756 438090 512778 438112
rect 512778 438090 512790 438112
rect 512856 438090 512868 438112
rect 512868 438090 512890 438112
rect 512956 438090 512958 438112
rect 512958 438090 512990 438112
rect 512756 438078 512790 438090
rect 512856 438078 512890 438090
rect 512956 438078 512990 438090
rect 513056 438078 513090 438112
rect 513156 438078 513190 438112
rect 513256 438090 513284 438112
rect 513284 438090 513290 438112
rect 513256 438078 513290 438090
rect 512756 438000 512778 438012
rect 512778 438000 512790 438012
rect 512856 438000 512868 438012
rect 512868 438000 512890 438012
rect 512956 438000 512958 438012
rect 512958 438000 512990 438012
rect 512756 437978 512790 438000
rect 512856 437978 512890 438000
rect 512956 437978 512990 438000
rect 513056 437978 513090 438012
rect 513156 437978 513190 438012
rect 513256 438000 513284 438012
rect 513284 438000 513290 438012
rect 513256 437978 513290 438000
rect 512756 437910 512778 437912
rect 512778 437910 512790 437912
rect 512856 437910 512868 437912
rect 512868 437910 512890 437912
rect 512956 437910 512958 437912
rect 512958 437910 512990 437912
rect 512756 437878 512790 437910
rect 512856 437878 512890 437910
rect 512956 437878 512990 437910
rect 513056 437878 513090 437912
rect 513156 437878 513190 437912
rect 513256 437910 513284 437912
rect 513284 437910 513290 437912
rect 513256 437878 513290 437910
rect 512756 437778 512790 437812
rect 512856 437778 512890 437812
rect 512956 437778 512990 437812
rect 513056 437778 513090 437812
rect 513156 437778 513190 437812
rect 513256 437778 513290 437812
rect 512756 437678 512790 437712
rect 512856 437678 512890 437712
rect 512956 437678 512990 437712
rect 513056 437678 513090 437712
rect 513156 437678 513190 437712
rect 513256 437678 513290 437712
rect 512756 437584 512790 437612
rect 512856 437584 512890 437612
rect 512956 437584 512990 437612
rect 512756 437578 512778 437584
rect 512778 437578 512790 437584
rect 512856 437578 512868 437584
rect 512868 437578 512890 437584
rect 512956 437578 512958 437584
rect 512958 437578 512990 437584
rect 513056 437578 513090 437612
rect 513156 437578 513190 437612
rect 513256 437584 513290 437612
rect 513256 437578 513284 437584
rect 513284 437578 513290 437584
rect 500418 437216 500518 437316
rect 500642 437216 500742 437316
rect 500866 437216 500966 437316
rect 501090 437216 501190 437316
rect 501314 437216 501368 437316
rect 501368 437216 501414 437316
rect 516208 438062 516605 438600
rect 522943 438062 523340 438600
rect 500418 436992 500518 437092
rect 500642 436992 500742 437092
rect 500866 436992 500966 437092
rect 501090 436992 501190 437092
rect 501314 436992 501368 437092
rect 501368 436992 501414 437092
rect 500418 436768 500518 436868
rect 500642 436768 500742 436868
rect 500866 436768 500966 436868
rect 501090 436768 501190 436868
rect 501314 436768 501368 436868
rect 501368 436768 501414 436868
rect 500418 436544 500518 436644
rect 500642 436544 500742 436644
rect 500866 436544 500966 436644
rect 501090 436544 501190 436644
rect 501314 436544 501368 436644
rect 501368 436544 501414 436644
rect 500418 436320 500518 436420
rect 500642 436320 500742 436420
rect 500866 436320 500966 436420
rect 501090 436320 501190 436420
rect 501314 436320 501368 436420
rect 501368 436320 501414 436420
rect 500418 436096 500518 436196
rect 500642 436096 500742 436196
rect 500866 436096 500966 436196
rect 501090 436096 501190 436196
rect 501314 436096 501368 436196
rect 501368 436096 501414 436196
rect 503740 436802 503762 436824
rect 503762 436802 503774 436824
rect 503840 436802 503852 436824
rect 503852 436802 503874 436824
rect 503940 436802 503942 436824
rect 503942 436802 503974 436824
rect 503740 436790 503774 436802
rect 503840 436790 503874 436802
rect 503940 436790 503974 436802
rect 504040 436790 504074 436824
rect 504140 436790 504174 436824
rect 504240 436802 504268 436824
rect 504268 436802 504274 436824
rect 504240 436790 504274 436802
rect 503740 436712 503762 436724
rect 503762 436712 503774 436724
rect 503840 436712 503852 436724
rect 503852 436712 503874 436724
rect 503940 436712 503942 436724
rect 503942 436712 503974 436724
rect 503740 436690 503774 436712
rect 503840 436690 503874 436712
rect 503940 436690 503974 436712
rect 504040 436690 504074 436724
rect 504140 436690 504174 436724
rect 504240 436712 504268 436724
rect 504268 436712 504274 436724
rect 504240 436690 504274 436712
rect 503740 436622 503762 436624
rect 503762 436622 503774 436624
rect 503840 436622 503852 436624
rect 503852 436622 503874 436624
rect 503940 436622 503942 436624
rect 503942 436622 503974 436624
rect 503740 436590 503774 436622
rect 503840 436590 503874 436622
rect 503940 436590 503974 436622
rect 504040 436590 504074 436624
rect 504140 436590 504174 436624
rect 504240 436622 504268 436624
rect 504268 436622 504274 436624
rect 504240 436590 504274 436622
rect 503740 436490 503774 436524
rect 503840 436490 503874 436524
rect 503940 436490 503974 436524
rect 504040 436490 504074 436524
rect 504140 436490 504174 436524
rect 504240 436490 504274 436524
rect 503740 436390 503774 436424
rect 503840 436390 503874 436424
rect 503940 436390 503974 436424
rect 504040 436390 504074 436424
rect 504140 436390 504174 436424
rect 504240 436390 504274 436424
rect 503740 436296 503774 436324
rect 503840 436296 503874 436324
rect 503940 436296 503974 436324
rect 503740 436290 503762 436296
rect 503762 436290 503774 436296
rect 503840 436290 503852 436296
rect 503852 436290 503874 436296
rect 503940 436290 503942 436296
rect 503942 436290 503974 436296
rect 504040 436290 504074 436324
rect 504140 436290 504174 436324
rect 504240 436296 504274 436324
rect 504240 436290 504268 436296
rect 504268 436290 504274 436296
rect 505028 436802 505050 436824
rect 505050 436802 505062 436824
rect 505128 436802 505140 436824
rect 505140 436802 505162 436824
rect 505228 436802 505230 436824
rect 505230 436802 505262 436824
rect 505028 436790 505062 436802
rect 505128 436790 505162 436802
rect 505228 436790 505262 436802
rect 505328 436790 505362 436824
rect 505428 436790 505462 436824
rect 505528 436802 505556 436824
rect 505556 436802 505562 436824
rect 505528 436790 505562 436802
rect 505028 436712 505050 436724
rect 505050 436712 505062 436724
rect 505128 436712 505140 436724
rect 505140 436712 505162 436724
rect 505228 436712 505230 436724
rect 505230 436712 505262 436724
rect 505028 436690 505062 436712
rect 505128 436690 505162 436712
rect 505228 436690 505262 436712
rect 505328 436690 505362 436724
rect 505428 436690 505462 436724
rect 505528 436712 505556 436724
rect 505556 436712 505562 436724
rect 505528 436690 505562 436712
rect 505028 436622 505050 436624
rect 505050 436622 505062 436624
rect 505128 436622 505140 436624
rect 505140 436622 505162 436624
rect 505228 436622 505230 436624
rect 505230 436622 505262 436624
rect 505028 436590 505062 436622
rect 505128 436590 505162 436622
rect 505228 436590 505262 436622
rect 505328 436590 505362 436624
rect 505428 436590 505462 436624
rect 505528 436622 505556 436624
rect 505556 436622 505562 436624
rect 505528 436590 505562 436622
rect 505028 436490 505062 436524
rect 505128 436490 505162 436524
rect 505228 436490 505262 436524
rect 505328 436490 505362 436524
rect 505428 436490 505462 436524
rect 505528 436490 505562 436524
rect 505028 436390 505062 436424
rect 505128 436390 505162 436424
rect 505228 436390 505262 436424
rect 505328 436390 505362 436424
rect 505428 436390 505462 436424
rect 505528 436390 505562 436424
rect 505028 436296 505062 436324
rect 505128 436296 505162 436324
rect 505228 436296 505262 436324
rect 505028 436290 505050 436296
rect 505050 436290 505062 436296
rect 505128 436290 505140 436296
rect 505140 436290 505162 436296
rect 505228 436290 505230 436296
rect 505230 436290 505262 436296
rect 505328 436290 505362 436324
rect 505428 436290 505462 436324
rect 505528 436296 505562 436324
rect 505528 436290 505556 436296
rect 505556 436290 505562 436296
rect 506316 436802 506338 436824
rect 506338 436802 506350 436824
rect 506416 436802 506428 436824
rect 506428 436802 506450 436824
rect 506516 436802 506518 436824
rect 506518 436802 506550 436824
rect 506316 436790 506350 436802
rect 506416 436790 506450 436802
rect 506516 436790 506550 436802
rect 506616 436790 506650 436824
rect 506716 436790 506750 436824
rect 506816 436802 506844 436824
rect 506844 436802 506850 436824
rect 506816 436790 506850 436802
rect 506316 436712 506338 436724
rect 506338 436712 506350 436724
rect 506416 436712 506428 436724
rect 506428 436712 506450 436724
rect 506516 436712 506518 436724
rect 506518 436712 506550 436724
rect 506316 436690 506350 436712
rect 506416 436690 506450 436712
rect 506516 436690 506550 436712
rect 506616 436690 506650 436724
rect 506716 436690 506750 436724
rect 506816 436712 506844 436724
rect 506844 436712 506850 436724
rect 506816 436690 506850 436712
rect 506316 436622 506338 436624
rect 506338 436622 506350 436624
rect 506416 436622 506428 436624
rect 506428 436622 506450 436624
rect 506516 436622 506518 436624
rect 506518 436622 506550 436624
rect 506316 436590 506350 436622
rect 506416 436590 506450 436622
rect 506516 436590 506550 436622
rect 506616 436590 506650 436624
rect 506716 436590 506750 436624
rect 506816 436622 506844 436624
rect 506844 436622 506850 436624
rect 506816 436590 506850 436622
rect 506316 436490 506350 436524
rect 506416 436490 506450 436524
rect 506516 436490 506550 436524
rect 506616 436490 506650 436524
rect 506716 436490 506750 436524
rect 506816 436490 506850 436524
rect 506316 436390 506350 436424
rect 506416 436390 506450 436424
rect 506516 436390 506550 436424
rect 506616 436390 506650 436424
rect 506716 436390 506750 436424
rect 506816 436390 506850 436424
rect 506316 436296 506350 436324
rect 506416 436296 506450 436324
rect 506516 436296 506550 436324
rect 506316 436290 506338 436296
rect 506338 436290 506350 436296
rect 506416 436290 506428 436296
rect 506428 436290 506450 436296
rect 506516 436290 506518 436296
rect 506518 436290 506550 436296
rect 506616 436290 506650 436324
rect 506716 436290 506750 436324
rect 506816 436296 506850 436324
rect 506816 436290 506844 436296
rect 506844 436290 506850 436296
rect 507604 436802 507626 436824
rect 507626 436802 507638 436824
rect 507704 436802 507716 436824
rect 507716 436802 507738 436824
rect 507804 436802 507806 436824
rect 507806 436802 507838 436824
rect 507604 436790 507638 436802
rect 507704 436790 507738 436802
rect 507804 436790 507838 436802
rect 507904 436790 507938 436824
rect 508004 436790 508038 436824
rect 508104 436802 508132 436824
rect 508132 436802 508138 436824
rect 508104 436790 508138 436802
rect 507604 436712 507626 436724
rect 507626 436712 507638 436724
rect 507704 436712 507716 436724
rect 507716 436712 507738 436724
rect 507804 436712 507806 436724
rect 507806 436712 507838 436724
rect 507604 436690 507638 436712
rect 507704 436690 507738 436712
rect 507804 436690 507838 436712
rect 507904 436690 507938 436724
rect 508004 436690 508038 436724
rect 508104 436712 508132 436724
rect 508132 436712 508138 436724
rect 508104 436690 508138 436712
rect 507604 436622 507626 436624
rect 507626 436622 507638 436624
rect 507704 436622 507716 436624
rect 507716 436622 507738 436624
rect 507804 436622 507806 436624
rect 507806 436622 507838 436624
rect 507604 436590 507638 436622
rect 507704 436590 507738 436622
rect 507804 436590 507838 436622
rect 507904 436590 507938 436624
rect 508004 436590 508038 436624
rect 508104 436622 508132 436624
rect 508132 436622 508138 436624
rect 508104 436590 508138 436622
rect 507604 436490 507638 436524
rect 507704 436490 507738 436524
rect 507804 436490 507838 436524
rect 507904 436490 507938 436524
rect 508004 436490 508038 436524
rect 508104 436490 508138 436524
rect 507604 436390 507638 436424
rect 507704 436390 507738 436424
rect 507804 436390 507838 436424
rect 507904 436390 507938 436424
rect 508004 436390 508038 436424
rect 508104 436390 508138 436424
rect 507604 436296 507638 436324
rect 507704 436296 507738 436324
rect 507804 436296 507838 436324
rect 507604 436290 507626 436296
rect 507626 436290 507638 436296
rect 507704 436290 507716 436296
rect 507716 436290 507738 436296
rect 507804 436290 507806 436296
rect 507806 436290 507838 436296
rect 507904 436290 507938 436324
rect 508004 436290 508038 436324
rect 508104 436296 508138 436324
rect 508104 436290 508132 436296
rect 508132 436290 508138 436296
rect 508892 436802 508914 436824
rect 508914 436802 508926 436824
rect 508992 436802 509004 436824
rect 509004 436802 509026 436824
rect 509092 436802 509094 436824
rect 509094 436802 509126 436824
rect 508892 436790 508926 436802
rect 508992 436790 509026 436802
rect 509092 436790 509126 436802
rect 509192 436790 509226 436824
rect 509292 436790 509326 436824
rect 509392 436802 509420 436824
rect 509420 436802 509426 436824
rect 509392 436790 509426 436802
rect 508892 436712 508914 436724
rect 508914 436712 508926 436724
rect 508992 436712 509004 436724
rect 509004 436712 509026 436724
rect 509092 436712 509094 436724
rect 509094 436712 509126 436724
rect 508892 436690 508926 436712
rect 508992 436690 509026 436712
rect 509092 436690 509126 436712
rect 509192 436690 509226 436724
rect 509292 436690 509326 436724
rect 509392 436712 509420 436724
rect 509420 436712 509426 436724
rect 509392 436690 509426 436712
rect 508892 436622 508914 436624
rect 508914 436622 508926 436624
rect 508992 436622 509004 436624
rect 509004 436622 509026 436624
rect 509092 436622 509094 436624
rect 509094 436622 509126 436624
rect 508892 436590 508926 436622
rect 508992 436590 509026 436622
rect 509092 436590 509126 436622
rect 509192 436590 509226 436624
rect 509292 436590 509326 436624
rect 509392 436622 509420 436624
rect 509420 436622 509426 436624
rect 509392 436590 509426 436622
rect 508892 436490 508926 436524
rect 508992 436490 509026 436524
rect 509092 436490 509126 436524
rect 509192 436490 509226 436524
rect 509292 436490 509326 436524
rect 509392 436490 509426 436524
rect 508892 436390 508926 436424
rect 508992 436390 509026 436424
rect 509092 436390 509126 436424
rect 509192 436390 509226 436424
rect 509292 436390 509326 436424
rect 509392 436390 509426 436424
rect 508892 436296 508926 436324
rect 508992 436296 509026 436324
rect 509092 436296 509126 436324
rect 508892 436290 508914 436296
rect 508914 436290 508926 436296
rect 508992 436290 509004 436296
rect 509004 436290 509026 436296
rect 509092 436290 509094 436296
rect 509094 436290 509126 436296
rect 509192 436290 509226 436324
rect 509292 436290 509326 436324
rect 509392 436296 509426 436324
rect 509392 436290 509420 436296
rect 509420 436290 509426 436296
rect 510180 436802 510202 436824
rect 510202 436802 510214 436824
rect 510280 436802 510292 436824
rect 510292 436802 510314 436824
rect 510380 436802 510382 436824
rect 510382 436802 510414 436824
rect 510180 436790 510214 436802
rect 510280 436790 510314 436802
rect 510380 436790 510414 436802
rect 510480 436790 510514 436824
rect 510580 436790 510614 436824
rect 510680 436802 510708 436824
rect 510708 436802 510714 436824
rect 510680 436790 510714 436802
rect 510180 436712 510202 436724
rect 510202 436712 510214 436724
rect 510280 436712 510292 436724
rect 510292 436712 510314 436724
rect 510380 436712 510382 436724
rect 510382 436712 510414 436724
rect 510180 436690 510214 436712
rect 510280 436690 510314 436712
rect 510380 436690 510414 436712
rect 510480 436690 510514 436724
rect 510580 436690 510614 436724
rect 510680 436712 510708 436724
rect 510708 436712 510714 436724
rect 510680 436690 510714 436712
rect 510180 436622 510202 436624
rect 510202 436622 510214 436624
rect 510280 436622 510292 436624
rect 510292 436622 510314 436624
rect 510380 436622 510382 436624
rect 510382 436622 510414 436624
rect 510180 436590 510214 436622
rect 510280 436590 510314 436622
rect 510380 436590 510414 436622
rect 510480 436590 510514 436624
rect 510580 436590 510614 436624
rect 510680 436622 510708 436624
rect 510708 436622 510714 436624
rect 510680 436590 510714 436622
rect 510180 436490 510214 436524
rect 510280 436490 510314 436524
rect 510380 436490 510414 436524
rect 510480 436490 510514 436524
rect 510580 436490 510614 436524
rect 510680 436490 510714 436524
rect 510180 436390 510214 436424
rect 510280 436390 510314 436424
rect 510380 436390 510414 436424
rect 510480 436390 510514 436424
rect 510580 436390 510614 436424
rect 510680 436390 510714 436424
rect 510180 436296 510214 436324
rect 510280 436296 510314 436324
rect 510380 436296 510414 436324
rect 510180 436290 510202 436296
rect 510202 436290 510214 436296
rect 510280 436290 510292 436296
rect 510292 436290 510314 436296
rect 510380 436290 510382 436296
rect 510382 436290 510414 436296
rect 510480 436290 510514 436324
rect 510580 436290 510614 436324
rect 510680 436296 510714 436324
rect 510680 436290 510708 436296
rect 510708 436290 510714 436296
rect 511468 436802 511490 436824
rect 511490 436802 511502 436824
rect 511568 436802 511580 436824
rect 511580 436802 511602 436824
rect 511668 436802 511670 436824
rect 511670 436802 511702 436824
rect 511468 436790 511502 436802
rect 511568 436790 511602 436802
rect 511668 436790 511702 436802
rect 511768 436790 511802 436824
rect 511868 436790 511902 436824
rect 511968 436802 511996 436824
rect 511996 436802 512002 436824
rect 511968 436790 512002 436802
rect 511468 436712 511490 436724
rect 511490 436712 511502 436724
rect 511568 436712 511580 436724
rect 511580 436712 511602 436724
rect 511668 436712 511670 436724
rect 511670 436712 511702 436724
rect 511468 436690 511502 436712
rect 511568 436690 511602 436712
rect 511668 436690 511702 436712
rect 511768 436690 511802 436724
rect 511868 436690 511902 436724
rect 511968 436712 511996 436724
rect 511996 436712 512002 436724
rect 511968 436690 512002 436712
rect 511468 436622 511490 436624
rect 511490 436622 511502 436624
rect 511568 436622 511580 436624
rect 511580 436622 511602 436624
rect 511668 436622 511670 436624
rect 511670 436622 511702 436624
rect 511468 436590 511502 436622
rect 511568 436590 511602 436622
rect 511668 436590 511702 436622
rect 511768 436590 511802 436624
rect 511868 436590 511902 436624
rect 511968 436622 511996 436624
rect 511996 436622 512002 436624
rect 511968 436590 512002 436622
rect 511468 436490 511502 436524
rect 511568 436490 511602 436524
rect 511668 436490 511702 436524
rect 511768 436490 511802 436524
rect 511868 436490 511902 436524
rect 511968 436490 512002 436524
rect 511468 436390 511502 436424
rect 511568 436390 511602 436424
rect 511668 436390 511702 436424
rect 511768 436390 511802 436424
rect 511868 436390 511902 436424
rect 511968 436390 512002 436424
rect 511468 436296 511502 436324
rect 511568 436296 511602 436324
rect 511668 436296 511702 436324
rect 511468 436290 511490 436296
rect 511490 436290 511502 436296
rect 511568 436290 511580 436296
rect 511580 436290 511602 436296
rect 511668 436290 511670 436296
rect 511670 436290 511702 436296
rect 511768 436290 511802 436324
rect 511868 436290 511902 436324
rect 511968 436296 512002 436324
rect 511968 436290 511996 436296
rect 511996 436290 512002 436296
rect 512756 436802 512778 436824
rect 512778 436802 512790 436824
rect 512856 436802 512868 436824
rect 512868 436802 512890 436824
rect 512956 436802 512958 436824
rect 512958 436802 512990 436824
rect 512756 436790 512790 436802
rect 512856 436790 512890 436802
rect 512956 436790 512990 436802
rect 513056 436790 513090 436824
rect 513156 436790 513190 436824
rect 513256 436802 513284 436824
rect 513284 436802 513290 436824
rect 513256 436790 513290 436802
rect 512756 436712 512778 436724
rect 512778 436712 512790 436724
rect 512856 436712 512868 436724
rect 512868 436712 512890 436724
rect 512956 436712 512958 436724
rect 512958 436712 512990 436724
rect 512756 436690 512790 436712
rect 512856 436690 512890 436712
rect 512956 436690 512990 436712
rect 513056 436690 513090 436724
rect 513156 436690 513190 436724
rect 513256 436712 513284 436724
rect 513284 436712 513290 436724
rect 513256 436690 513290 436712
rect 512756 436622 512778 436624
rect 512778 436622 512790 436624
rect 512856 436622 512868 436624
rect 512868 436622 512890 436624
rect 512956 436622 512958 436624
rect 512958 436622 512990 436624
rect 512756 436590 512790 436622
rect 512856 436590 512890 436622
rect 512956 436590 512990 436622
rect 513056 436590 513090 436624
rect 513156 436590 513190 436624
rect 513256 436622 513284 436624
rect 513284 436622 513290 436624
rect 513256 436590 513290 436622
rect 512756 436490 512790 436524
rect 512856 436490 512890 436524
rect 512956 436490 512990 436524
rect 513056 436490 513090 436524
rect 513156 436490 513190 436524
rect 513256 436490 513290 436524
rect 512756 436390 512790 436424
rect 512856 436390 512890 436424
rect 512956 436390 512990 436424
rect 513056 436390 513090 436424
rect 513156 436390 513190 436424
rect 513256 436390 513290 436424
rect 512756 436296 512790 436324
rect 512856 436296 512890 436324
rect 512956 436296 512990 436324
rect 512756 436290 512778 436296
rect 512778 436290 512790 436296
rect 512856 436290 512868 436296
rect 512868 436290 512890 436296
rect 512956 436290 512958 436296
rect 512958 436290 512990 436296
rect 513056 436290 513090 436324
rect 513156 436290 513190 436324
rect 513256 436296 513290 436324
rect 513256 436290 513284 436296
rect 513284 436290 513290 436296
rect 500418 435872 500518 435972
rect 500642 435872 500742 435972
rect 500866 435872 500966 435972
rect 501090 435872 501190 435972
rect 501314 435872 501368 435972
rect 501368 435872 501414 435972
rect 500418 435648 500518 435748
rect 500642 435648 500742 435748
rect 500866 435648 500966 435748
rect 501090 435648 501190 435748
rect 501314 435648 501368 435748
rect 501368 435648 501414 435748
rect 500418 435424 500518 435524
rect 500642 435424 500742 435524
rect 500866 435424 500966 435524
rect 501090 435424 501190 435524
rect 501314 435424 501368 435524
rect 501368 435424 501414 435524
rect 500418 435200 500518 435300
rect 500642 435200 500742 435300
rect 500866 435200 500966 435300
rect 501090 435200 501190 435300
rect 501314 435200 501368 435300
rect 501368 435200 501414 435300
rect 500418 434976 500518 435076
rect 500642 434976 500742 435076
rect 500866 434976 500966 435076
rect 501090 434976 501190 435076
rect 501314 434976 501368 435076
rect 501368 434976 501414 435076
rect 503740 435514 503762 435536
rect 503762 435514 503774 435536
rect 503840 435514 503852 435536
rect 503852 435514 503874 435536
rect 503940 435514 503942 435536
rect 503942 435514 503974 435536
rect 503740 435502 503774 435514
rect 503840 435502 503874 435514
rect 503940 435502 503974 435514
rect 504040 435502 504074 435536
rect 504140 435502 504174 435536
rect 504240 435514 504268 435536
rect 504268 435514 504274 435536
rect 504240 435502 504274 435514
rect 503740 435424 503762 435436
rect 503762 435424 503774 435436
rect 503840 435424 503852 435436
rect 503852 435424 503874 435436
rect 503940 435424 503942 435436
rect 503942 435424 503974 435436
rect 503740 435402 503774 435424
rect 503840 435402 503874 435424
rect 503940 435402 503974 435424
rect 504040 435402 504074 435436
rect 504140 435402 504174 435436
rect 504240 435424 504268 435436
rect 504268 435424 504274 435436
rect 504240 435402 504274 435424
rect 503740 435334 503762 435336
rect 503762 435334 503774 435336
rect 503840 435334 503852 435336
rect 503852 435334 503874 435336
rect 503940 435334 503942 435336
rect 503942 435334 503974 435336
rect 503740 435302 503774 435334
rect 503840 435302 503874 435334
rect 503940 435302 503974 435334
rect 504040 435302 504074 435336
rect 504140 435302 504174 435336
rect 504240 435334 504268 435336
rect 504268 435334 504274 435336
rect 504240 435302 504274 435334
rect 503740 435202 503774 435236
rect 503840 435202 503874 435236
rect 503940 435202 503974 435236
rect 504040 435202 504074 435236
rect 504140 435202 504174 435236
rect 504240 435202 504274 435236
rect 503740 435102 503774 435136
rect 503840 435102 503874 435136
rect 503940 435102 503974 435136
rect 504040 435102 504074 435136
rect 504140 435102 504174 435136
rect 504240 435102 504274 435136
rect 503740 435008 503774 435036
rect 503840 435008 503874 435036
rect 503940 435008 503974 435036
rect 503740 435002 503762 435008
rect 503762 435002 503774 435008
rect 503840 435002 503852 435008
rect 503852 435002 503874 435008
rect 503940 435002 503942 435008
rect 503942 435002 503974 435008
rect 504040 435002 504074 435036
rect 504140 435002 504174 435036
rect 504240 435008 504274 435036
rect 504240 435002 504268 435008
rect 504268 435002 504274 435008
rect 500418 434752 500518 434852
rect 500642 434752 500742 434852
rect 500866 434752 500966 434852
rect 501090 434752 501190 434852
rect 501314 434752 501368 434852
rect 501368 434752 501414 434852
rect 505028 435514 505050 435536
rect 505050 435514 505062 435536
rect 505128 435514 505140 435536
rect 505140 435514 505162 435536
rect 505228 435514 505230 435536
rect 505230 435514 505262 435536
rect 505028 435502 505062 435514
rect 505128 435502 505162 435514
rect 505228 435502 505262 435514
rect 505328 435502 505362 435536
rect 505428 435502 505462 435536
rect 505528 435514 505556 435536
rect 505556 435514 505562 435536
rect 505528 435502 505562 435514
rect 505028 435424 505050 435436
rect 505050 435424 505062 435436
rect 505128 435424 505140 435436
rect 505140 435424 505162 435436
rect 505228 435424 505230 435436
rect 505230 435424 505262 435436
rect 505028 435402 505062 435424
rect 505128 435402 505162 435424
rect 505228 435402 505262 435424
rect 505328 435402 505362 435436
rect 505428 435402 505462 435436
rect 505528 435424 505556 435436
rect 505556 435424 505562 435436
rect 505528 435402 505562 435424
rect 505028 435334 505050 435336
rect 505050 435334 505062 435336
rect 505128 435334 505140 435336
rect 505140 435334 505162 435336
rect 505228 435334 505230 435336
rect 505230 435334 505262 435336
rect 505028 435302 505062 435334
rect 505128 435302 505162 435334
rect 505228 435302 505262 435334
rect 505328 435302 505362 435336
rect 505428 435302 505462 435336
rect 505528 435334 505556 435336
rect 505556 435334 505562 435336
rect 505528 435302 505562 435334
rect 505028 435202 505062 435236
rect 505128 435202 505162 435236
rect 505228 435202 505262 435236
rect 505328 435202 505362 435236
rect 505428 435202 505462 435236
rect 505528 435202 505562 435236
rect 505028 435102 505062 435136
rect 505128 435102 505162 435136
rect 505228 435102 505262 435136
rect 505328 435102 505362 435136
rect 505428 435102 505462 435136
rect 505528 435102 505562 435136
rect 505028 435008 505062 435036
rect 505128 435008 505162 435036
rect 505228 435008 505262 435036
rect 505028 435002 505050 435008
rect 505050 435002 505062 435008
rect 505128 435002 505140 435008
rect 505140 435002 505162 435008
rect 505228 435002 505230 435008
rect 505230 435002 505262 435008
rect 505328 435002 505362 435036
rect 505428 435002 505462 435036
rect 505528 435008 505562 435036
rect 505528 435002 505556 435008
rect 505556 435002 505562 435008
rect 506316 435514 506338 435536
rect 506338 435514 506350 435536
rect 506416 435514 506428 435536
rect 506428 435514 506450 435536
rect 506516 435514 506518 435536
rect 506518 435514 506550 435536
rect 506316 435502 506350 435514
rect 506416 435502 506450 435514
rect 506516 435502 506550 435514
rect 506616 435502 506650 435536
rect 506716 435502 506750 435536
rect 506816 435514 506844 435536
rect 506844 435514 506850 435536
rect 506816 435502 506850 435514
rect 506316 435424 506338 435436
rect 506338 435424 506350 435436
rect 506416 435424 506428 435436
rect 506428 435424 506450 435436
rect 506516 435424 506518 435436
rect 506518 435424 506550 435436
rect 506316 435402 506350 435424
rect 506416 435402 506450 435424
rect 506516 435402 506550 435424
rect 506616 435402 506650 435436
rect 506716 435402 506750 435436
rect 506816 435424 506844 435436
rect 506844 435424 506850 435436
rect 506816 435402 506850 435424
rect 506316 435334 506338 435336
rect 506338 435334 506350 435336
rect 506416 435334 506428 435336
rect 506428 435334 506450 435336
rect 506516 435334 506518 435336
rect 506518 435334 506550 435336
rect 506316 435302 506350 435334
rect 506416 435302 506450 435334
rect 506516 435302 506550 435334
rect 506616 435302 506650 435336
rect 506716 435302 506750 435336
rect 506816 435334 506844 435336
rect 506844 435334 506850 435336
rect 506816 435302 506850 435334
rect 506316 435202 506350 435236
rect 506416 435202 506450 435236
rect 506516 435202 506550 435236
rect 506616 435202 506650 435236
rect 506716 435202 506750 435236
rect 506816 435202 506850 435236
rect 506316 435102 506350 435136
rect 506416 435102 506450 435136
rect 506516 435102 506550 435136
rect 506616 435102 506650 435136
rect 506716 435102 506750 435136
rect 506816 435102 506850 435136
rect 506316 435008 506350 435036
rect 506416 435008 506450 435036
rect 506516 435008 506550 435036
rect 506316 435002 506338 435008
rect 506338 435002 506350 435008
rect 506416 435002 506428 435008
rect 506428 435002 506450 435008
rect 506516 435002 506518 435008
rect 506518 435002 506550 435008
rect 506616 435002 506650 435036
rect 506716 435002 506750 435036
rect 506816 435008 506850 435036
rect 506816 435002 506844 435008
rect 506844 435002 506850 435008
rect 507604 435514 507626 435536
rect 507626 435514 507638 435536
rect 507704 435514 507716 435536
rect 507716 435514 507738 435536
rect 507804 435514 507806 435536
rect 507806 435514 507838 435536
rect 507604 435502 507638 435514
rect 507704 435502 507738 435514
rect 507804 435502 507838 435514
rect 507904 435502 507938 435536
rect 508004 435502 508038 435536
rect 508104 435514 508132 435536
rect 508132 435514 508138 435536
rect 508104 435502 508138 435514
rect 507604 435424 507626 435436
rect 507626 435424 507638 435436
rect 507704 435424 507716 435436
rect 507716 435424 507738 435436
rect 507804 435424 507806 435436
rect 507806 435424 507838 435436
rect 507604 435402 507638 435424
rect 507704 435402 507738 435424
rect 507804 435402 507838 435424
rect 507904 435402 507938 435436
rect 508004 435402 508038 435436
rect 508104 435424 508132 435436
rect 508132 435424 508138 435436
rect 508104 435402 508138 435424
rect 507604 435334 507626 435336
rect 507626 435334 507638 435336
rect 507704 435334 507716 435336
rect 507716 435334 507738 435336
rect 507804 435334 507806 435336
rect 507806 435334 507838 435336
rect 507604 435302 507638 435334
rect 507704 435302 507738 435334
rect 507804 435302 507838 435334
rect 507904 435302 507938 435336
rect 508004 435302 508038 435336
rect 508104 435334 508132 435336
rect 508132 435334 508138 435336
rect 508104 435302 508138 435334
rect 507604 435202 507638 435236
rect 507704 435202 507738 435236
rect 507804 435202 507838 435236
rect 507904 435202 507938 435236
rect 508004 435202 508038 435236
rect 508104 435202 508138 435236
rect 507604 435102 507638 435136
rect 507704 435102 507738 435136
rect 507804 435102 507838 435136
rect 507904 435102 507938 435136
rect 508004 435102 508038 435136
rect 508104 435102 508138 435136
rect 507604 435008 507638 435036
rect 507704 435008 507738 435036
rect 507804 435008 507838 435036
rect 507604 435002 507626 435008
rect 507626 435002 507638 435008
rect 507704 435002 507716 435008
rect 507716 435002 507738 435008
rect 507804 435002 507806 435008
rect 507806 435002 507838 435008
rect 507904 435002 507938 435036
rect 508004 435002 508038 435036
rect 508104 435008 508138 435036
rect 508104 435002 508132 435008
rect 508132 435002 508138 435008
rect 508892 435514 508914 435536
rect 508914 435514 508926 435536
rect 508992 435514 509004 435536
rect 509004 435514 509026 435536
rect 509092 435514 509094 435536
rect 509094 435514 509126 435536
rect 508892 435502 508926 435514
rect 508992 435502 509026 435514
rect 509092 435502 509126 435514
rect 509192 435502 509226 435536
rect 509292 435502 509326 435536
rect 509392 435514 509420 435536
rect 509420 435514 509426 435536
rect 509392 435502 509426 435514
rect 508892 435424 508914 435436
rect 508914 435424 508926 435436
rect 508992 435424 509004 435436
rect 509004 435424 509026 435436
rect 509092 435424 509094 435436
rect 509094 435424 509126 435436
rect 508892 435402 508926 435424
rect 508992 435402 509026 435424
rect 509092 435402 509126 435424
rect 509192 435402 509226 435436
rect 509292 435402 509326 435436
rect 509392 435424 509420 435436
rect 509420 435424 509426 435436
rect 509392 435402 509426 435424
rect 508892 435334 508914 435336
rect 508914 435334 508926 435336
rect 508992 435334 509004 435336
rect 509004 435334 509026 435336
rect 509092 435334 509094 435336
rect 509094 435334 509126 435336
rect 508892 435302 508926 435334
rect 508992 435302 509026 435334
rect 509092 435302 509126 435334
rect 509192 435302 509226 435336
rect 509292 435302 509326 435336
rect 509392 435334 509420 435336
rect 509420 435334 509426 435336
rect 509392 435302 509426 435334
rect 508892 435202 508926 435236
rect 508992 435202 509026 435236
rect 509092 435202 509126 435236
rect 509192 435202 509226 435236
rect 509292 435202 509326 435236
rect 509392 435202 509426 435236
rect 508892 435102 508926 435136
rect 508992 435102 509026 435136
rect 509092 435102 509126 435136
rect 509192 435102 509226 435136
rect 509292 435102 509326 435136
rect 509392 435102 509426 435136
rect 508892 435008 508926 435036
rect 508992 435008 509026 435036
rect 509092 435008 509126 435036
rect 508892 435002 508914 435008
rect 508914 435002 508926 435008
rect 508992 435002 509004 435008
rect 509004 435002 509026 435008
rect 509092 435002 509094 435008
rect 509094 435002 509126 435008
rect 509192 435002 509226 435036
rect 509292 435002 509326 435036
rect 509392 435008 509426 435036
rect 509392 435002 509420 435008
rect 509420 435002 509426 435008
rect 510180 435514 510202 435536
rect 510202 435514 510214 435536
rect 510280 435514 510292 435536
rect 510292 435514 510314 435536
rect 510380 435514 510382 435536
rect 510382 435514 510414 435536
rect 510180 435502 510214 435514
rect 510280 435502 510314 435514
rect 510380 435502 510414 435514
rect 510480 435502 510514 435536
rect 510580 435502 510614 435536
rect 510680 435514 510708 435536
rect 510708 435514 510714 435536
rect 510680 435502 510714 435514
rect 510180 435424 510202 435436
rect 510202 435424 510214 435436
rect 510280 435424 510292 435436
rect 510292 435424 510314 435436
rect 510380 435424 510382 435436
rect 510382 435424 510414 435436
rect 510180 435402 510214 435424
rect 510280 435402 510314 435424
rect 510380 435402 510414 435424
rect 510480 435402 510514 435436
rect 510580 435402 510614 435436
rect 510680 435424 510708 435436
rect 510708 435424 510714 435436
rect 510680 435402 510714 435424
rect 510180 435334 510202 435336
rect 510202 435334 510214 435336
rect 510280 435334 510292 435336
rect 510292 435334 510314 435336
rect 510380 435334 510382 435336
rect 510382 435334 510414 435336
rect 510180 435302 510214 435334
rect 510280 435302 510314 435334
rect 510380 435302 510414 435334
rect 510480 435302 510514 435336
rect 510580 435302 510614 435336
rect 510680 435334 510708 435336
rect 510708 435334 510714 435336
rect 510680 435302 510714 435334
rect 510180 435202 510214 435236
rect 510280 435202 510314 435236
rect 510380 435202 510414 435236
rect 510480 435202 510514 435236
rect 510580 435202 510614 435236
rect 510680 435202 510714 435236
rect 510180 435102 510214 435136
rect 510280 435102 510314 435136
rect 510380 435102 510414 435136
rect 510480 435102 510514 435136
rect 510580 435102 510614 435136
rect 510680 435102 510714 435136
rect 510180 435008 510214 435036
rect 510280 435008 510314 435036
rect 510380 435008 510414 435036
rect 510180 435002 510202 435008
rect 510202 435002 510214 435008
rect 510280 435002 510292 435008
rect 510292 435002 510314 435008
rect 510380 435002 510382 435008
rect 510382 435002 510414 435008
rect 510480 435002 510514 435036
rect 510580 435002 510614 435036
rect 510680 435008 510714 435036
rect 510680 435002 510708 435008
rect 510708 435002 510714 435008
rect 511468 435514 511490 435536
rect 511490 435514 511502 435536
rect 511568 435514 511580 435536
rect 511580 435514 511602 435536
rect 511668 435514 511670 435536
rect 511670 435514 511702 435536
rect 511468 435502 511502 435514
rect 511568 435502 511602 435514
rect 511668 435502 511702 435514
rect 511768 435502 511802 435536
rect 511868 435502 511902 435536
rect 511968 435514 511996 435536
rect 511996 435514 512002 435536
rect 511968 435502 512002 435514
rect 511468 435424 511490 435436
rect 511490 435424 511502 435436
rect 511568 435424 511580 435436
rect 511580 435424 511602 435436
rect 511668 435424 511670 435436
rect 511670 435424 511702 435436
rect 511468 435402 511502 435424
rect 511568 435402 511602 435424
rect 511668 435402 511702 435424
rect 511768 435402 511802 435436
rect 511868 435402 511902 435436
rect 511968 435424 511996 435436
rect 511996 435424 512002 435436
rect 511968 435402 512002 435424
rect 511468 435334 511490 435336
rect 511490 435334 511502 435336
rect 511568 435334 511580 435336
rect 511580 435334 511602 435336
rect 511668 435334 511670 435336
rect 511670 435334 511702 435336
rect 511468 435302 511502 435334
rect 511568 435302 511602 435334
rect 511668 435302 511702 435334
rect 511768 435302 511802 435336
rect 511868 435302 511902 435336
rect 511968 435334 511996 435336
rect 511996 435334 512002 435336
rect 511968 435302 512002 435334
rect 511468 435202 511502 435236
rect 511568 435202 511602 435236
rect 511668 435202 511702 435236
rect 511768 435202 511802 435236
rect 511868 435202 511902 435236
rect 511968 435202 512002 435236
rect 511468 435102 511502 435136
rect 511568 435102 511602 435136
rect 511668 435102 511702 435136
rect 511768 435102 511802 435136
rect 511868 435102 511902 435136
rect 511968 435102 512002 435136
rect 511468 435008 511502 435036
rect 511568 435008 511602 435036
rect 511668 435008 511702 435036
rect 511468 435002 511490 435008
rect 511490 435002 511502 435008
rect 511568 435002 511580 435008
rect 511580 435002 511602 435008
rect 511668 435002 511670 435008
rect 511670 435002 511702 435008
rect 511768 435002 511802 435036
rect 511868 435002 511902 435036
rect 511968 435008 512002 435036
rect 511968 435002 511996 435008
rect 511996 435002 512002 435008
rect 512756 435514 512778 435536
rect 512778 435514 512790 435536
rect 512856 435514 512868 435536
rect 512868 435514 512890 435536
rect 512956 435514 512958 435536
rect 512958 435514 512990 435536
rect 512756 435502 512790 435514
rect 512856 435502 512890 435514
rect 512956 435502 512990 435514
rect 513056 435502 513090 435536
rect 513156 435502 513190 435536
rect 513256 435514 513284 435536
rect 513284 435514 513290 435536
rect 513256 435502 513290 435514
rect 512756 435424 512778 435436
rect 512778 435424 512790 435436
rect 512856 435424 512868 435436
rect 512868 435424 512890 435436
rect 512956 435424 512958 435436
rect 512958 435424 512990 435436
rect 512756 435402 512790 435424
rect 512856 435402 512890 435424
rect 512956 435402 512990 435424
rect 513056 435402 513090 435436
rect 513156 435402 513190 435436
rect 513256 435424 513284 435436
rect 513284 435424 513290 435436
rect 513256 435402 513290 435424
rect 512756 435334 512778 435336
rect 512778 435334 512790 435336
rect 512856 435334 512868 435336
rect 512868 435334 512890 435336
rect 512956 435334 512958 435336
rect 512958 435334 512990 435336
rect 512756 435302 512790 435334
rect 512856 435302 512890 435334
rect 512956 435302 512990 435334
rect 513056 435302 513090 435336
rect 513156 435302 513190 435336
rect 513256 435334 513284 435336
rect 513284 435334 513290 435336
rect 513256 435302 513290 435334
rect 512756 435202 512790 435236
rect 512856 435202 512890 435236
rect 512956 435202 512990 435236
rect 513056 435202 513090 435236
rect 513156 435202 513190 435236
rect 513256 435202 513290 435236
rect 512756 435102 512790 435136
rect 512856 435102 512890 435136
rect 512956 435102 512990 435136
rect 513056 435102 513090 435136
rect 513156 435102 513190 435136
rect 513256 435102 513290 435136
rect 512756 435008 512790 435036
rect 512856 435008 512890 435036
rect 512956 435008 512990 435036
rect 512756 435002 512778 435008
rect 512778 435002 512790 435008
rect 512856 435002 512868 435008
rect 512868 435002 512890 435008
rect 512956 435002 512958 435008
rect 512958 435002 512990 435008
rect 513056 435002 513090 435036
rect 513156 435002 513190 435036
rect 513256 435008 513290 435036
rect 513256 435002 513284 435008
rect 513284 435002 513290 435008
rect 500418 434528 500518 434628
rect 500642 434528 500742 434628
rect 500866 434528 500966 434628
rect 501090 434528 501190 434628
rect 501314 434528 501368 434628
rect 501368 434528 501414 434628
rect 500418 434304 500518 434404
rect 500642 434304 500742 434404
rect 500866 434304 500966 434404
rect 501090 434304 501190 434404
rect 501314 434304 501368 434404
rect 501368 434304 501414 434404
rect 500418 434080 500518 434180
rect 500642 434080 500742 434180
rect 500866 434080 500966 434180
rect 501090 434080 501190 434180
rect 501314 434080 501368 434180
rect 501368 434080 501414 434180
rect 500418 433856 500518 433956
rect 500642 433856 500742 433956
rect 500866 433856 500966 433956
rect 501090 433856 501190 433956
rect 501314 433856 501368 433956
rect 501368 433856 501414 433956
rect 500418 433632 500518 433732
rect 500642 433632 500742 433732
rect 500866 433632 500966 433732
rect 501090 433632 501190 433732
rect 501314 433632 501368 433732
rect 501368 433632 501414 433732
rect 503740 434226 503762 434248
rect 503762 434226 503774 434248
rect 503840 434226 503852 434248
rect 503852 434226 503874 434248
rect 503940 434226 503942 434248
rect 503942 434226 503974 434248
rect 503740 434214 503774 434226
rect 503840 434214 503874 434226
rect 503940 434214 503974 434226
rect 504040 434214 504074 434248
rect 504140 434214 504174 434248
rect 504240 434226 504268 434248
rect 504268 434226 504274 434248
rect 504240 434214 504274 434226
rect 503740 434136 503762 434148
rect 503762 434136 503774 434148
rect 503840 434136 503852 434148
rect 503852 434136 503874 434148
rect 503940 434136 503942 434148
rect 503942 434136 503974 434148
rect 503740 434114 503774 434136
rect 503840 434114 503874 434136
rect 503940 434114 503974 434136
rect 504040 434114 504074 434148
rect 504140 434114 504174 434148
rect 504240 434136 504268 434148
rect 504268 434136 504274 434148
rect 504240 434114 504274 434136
rect 503740 434046 503762 434048
rect 503762 434046 503774 434048
rect 503840 434046 503852 434048
rect 503852 434046 503874 434048
rect 503940 434046 503942 434048
rect 503942 434046 503974 434048
rect 503740 434014 503774 434046
rect 503840 434014 503874 434046
rect 503940 434014 503974 434046
rect 504040 434014 504074 434048
rect 504140 434014 504174 434048
rect 504240 434046 504268 434048
rect 504268 434046 504274 434048
rect 504240 434014 504274 434046
rect 503740 433914 503774 433948
rect 503840 433914 503874 433948
rect 503940 433914 503974 433948
rect 504040 433914 504074 433948
rect 504140 433914 504174 433948
rect 504240 433914 504274 433948
rect 503740 433814 503774 433848
rect 503840 433814 503874 433848
rect 503940 433814 503974 433848
rect 504040 433814 504074 433848
rect 504140 433814 504174 433848
rect 504240 433814 504274 433848
rect 503740 433720 503774 433748
rect 503840 433720 503874 433748
rect 503940 433720 503974 433748
rect 503740 433714 503762 433720
rect 503762 433714 503774 433720
rect 503840 433714 503852 433720
rect 503852 433714 503874 433720
rect 503940 433714 503942 433720
rect 503942 433714 503974 433720
rect 504040 433714 504074 433748
rect 504140 433714 504174 433748
rect 504240 433720 504274 433748
rect 504240 433714 504268 433720
rect 504268 433714 504274 433720
rect 505028 434226 505050 434248
rect 505050 434226 505062 434248
rect 505128 434226 505140 434248
rect 505140 434226 505162 434248
rect 505228 434226 505230 434248
rect 505230 434226 505262 434248
rect 505028 434214 505062 434226
rect 505128 434214 505162 434226
rect 505228 434214 505262 434226
rect 505328 434214 505362 434248
rect 505428 434214 505462 434248
rect 505528 434226 505556 434248
rect 505556 434226 505562 434248
rect 505528 434214 505562 434226
rect 505028 434136 505050 434148
rect 505050 434136 505062 434148
rect 505128 434136 505140 434148
rect 505140 434136 505162 434148
rect 505228 434136 505230 434148
rect 505230 434136 505262 434148
rect 505028 434114 505062 434136
rect 505128 434114 505162 434136
rect 505228 434114 505262 434136
rect 505328 434114 505362 434148
rect 505428 434114 505462 434148
rect 505528 434136 505556 434148
rect 505556 434136 505562 434148
rect 505528 434114 505562 434136
rect 505028 434046 505050 434048
rect 505050 434046 505062 434048
rect 505128 434046 505140 434048
rect 505140 434046 505162 434048
rect 505228 434046 505230 434048
rect 505230 434046 505262 434048
rect 505028 434014 505062 434046
rect 505128 434014 505162 434046
rect 505228 434014 505262 434046
rect 505328 434014 505362 434048
rect 505428 434014 505462 434048
rect 505528 434046 505556 434048
rect 505556 434046 505562 434048
rect 505528 434014 505562 434046
rect 505028 433914 505062 433948
rect 505128 433914 505162 433948
rect 505228 433914 505262 433948
rect 505328 433914 505362 433948
rect 505428 433914 505462 433948
rect 505528 433914 505562 433948
rect 505028 433814 505062 433848
rect 505128 433814 505162 433848
rect 505228 433814 505262 433848
rect 505328 433814 505362 433848
rect 505428 433814 505462 433848
rect 505528 433814 505562 433848
rect 505028 433720 505062 433748
rect 505128 433720 505162 433748
rect 505228 433720 505262 433748
rect 505028 433714 505050 433720
rect 505050 433714 505062 433720
rect 505128 433714 505140 433720
rect 505140 433714 505162 433720
rect 505228 433714 505230 433720
rect 505230 433714 505262 433720
rect 505328 433714 505362 433748
rect 505428 433714 505462 433748
rect 505528 433720 505562 433748
rect 505528 433714 505556 433720
rect 505556 433714 505562 433720
rect 506316 434226 506338 434248
rect 506338 434226 506350 434248
rect 506416 434226 506428 434248
rect 506428 434226 506450 434248
rect 506516 434226 506518 434248
rect 506518 434226 506550 434248
rect 506316 434214 506350 434226
rect 506416 434214 506450 434226
rect 506516 434214 506550 434226
rect 506616 434214 506650 434248
rect 506716 434214 506750 434248
rect 506816 434226 506844 434248
rect 506844 434226 506850 434248
rect 506816 434214 506850 434226
rect 506316 434136 506338 434148
rect 506338 434136 506350 434148
rect 506416 434136 506428 434148
rect 506428 434136 506450 434148
rect 506516 434136 506518 434148
rect 506518 434136 506550 434148
rect 506316 434114 506350 434136
rect 506416 434114 506450 434136
rect 506516 434114 506550 434136
rect 506616 434114 506650 434148
rect 506716 434114 506750 434148
rect 506816 434136 506844 434148
rect 506844 434136 506850 434148
rect 506816 434114 506850 434136
rect 506316 434046 506338 434048
rect 506338 434046 506350 434048
rect 506416 434046 506428 434048
rect 506428 434046 506450 434048
rect 506516 434046 506518 434048
rect 506518 434046 506550 434048
rect 506316 434014 506350 434046
rect 506416 434014 506450 434046
rect 506516 434014 506550 434046
rect 506616 434014 506650 434048
rect 506716 434014 506750 434048
rect 506816 434046 506844 434048
rect 506844 434046 506850 434048
rect 506816 434014 506850 434046
rect 506316 433914 506350 433948
rect 506416 433914 506450 433948
rect 506516 433914 506550 433948
rect 506616 433914 506650 433948
rect 506716 433914 506750 433948
rect 506816 433914 506850 433948
rect 506316 433814 506350 433848
rect 506416 433814 506450 433848
rect 506516 433814 506550 433848
rect 506616 433814 506650 433848
rect 506716 433814 506750 433848
rect 506816 433814 506850 433848
rect 506316 433720 506350 433748
rect 506416 433720 506450 433748
rect 506516 433720 506550 433748
rect 506316 433714 506338 433720
rect 506338 433714 506350 433720
rect 506416 433714 506428 433720
rect 506428 433714 506450 433720
rect 506516 433714 506518 433720
rect 506518 433714 506550 433720
rect 506616 433714 506650 433748
rect 506716 433714 506750 433748
rect 506816 433720 506850 433748
rect 506816 433714 506844 433720
rect 506844 433714 506850 433720
rect 507604 434226 507626 434248
rect 507626 434226 507638 434248
rect 507704 434226 507716 434248
rect 507716 434226 507738 434248
rect 507804 434226 507806 434248
rect 507806 434226 507838 434248
rect 507604 434214 507638 434226
rect 507704 434214 507738 434226
rect 507804 434214 507838 434226
rect 507904 434214 507938 434248
rect 508004 434214 508038 434248
rect 508104 434226 508132 434248
rect 508132 434226 508138 434248
rect 508104 434214 508138 434226
rect 507604 434136 507626 434148
rect 507626 434136 507638 434148
rect 507704 434136 507716 434148
rect 507716 434136 507738 434148
rect 507804 434136 507806 434148
rect 507806 434136 507838 434148
rect 507604 434114 507638 434136
rect 507704 434114 507738 434136
rect 507804 434114 507838 434136
rect 507904 434114 507938 434148
rect 508004 434114 508038 434148
rect 508104 434136 508132 434148
rect 508132 434136 508138 434148
rect 508104 434114 508138 434136
rect 507604 434046 507626 434048
rect 507626 434046 507638 434048
rect 507704 434046 507716 434048
rect 507716 434046 507738 434048
rect 507804 434046 507806 434048
rect 507806 434046 507838 434048
rect 507604 434014 507638 434046
rect 507704 434014 507738 434046
rect 507804 434014 507838 434046
rect 507904 434014 507938 434048
rect 508004 434014 508038 434048
rect 508104 434046 508132 434048
rect 508132 434046 508138 434048
rect 508104 434014 508138 434046
rect 507604 433914 507638 433948
rect 507704 433914 507738 433948
rect 507804 433914 507838 433948
rect 507904 433914 507938 433948
rect 508004 433914 508038 433948
rect 508104 433914 508138 433948
rect 507604 433814 507638 433848
rect 507704 433814 507738 433848
rect 507804 433814 507838 433848
rect 507904 433814 507938 433848
rect 508004 433814 508038 433848
rect 508104 433814 508138 433848
rect 507604 433720 507638 433748
rect 507704 433720 507738 433748
rect 507804 433720 507838 433748
rect 507604 433714 507626 433720
rect 507626 433714 507638 433720
rect 507704 433714 507716 433720
rect 507716 433714 507738 433720
rect 507804 433714 507806 433720
rect 507806 433714 507838 433720
rect 507904 433714 507938 433748
rect 508004 433714 508038 433748
rect 508104 433720 508138 433748
rect 508104 433714 508132 433720
rect 508132 433714 508138 433720
rect 508892 434226 508914 434248
rect 508914 434226 508926 434248
rect 508992 434226 509004 434248
rect 509004 434226 509026 434248
rect 509092 434226 509094 434248
rect 509094 434226 509126 434248
rect 508892 434214 508926 434226
rect 508992 434214 509026 434226
rect 509092 434214 509126 434226
rect 509192 434214 509226 434248
rect 509292 434214 509326 434248
rect 509392 434226 509420 434248
rect 509420 434226 509426 434248
rect 509392 434214 509426 434226
rect 508892 434136 508914 434148
rect 508914 434136 508926 434148
rect 508992 434136 509004 434148
rect 509004 434136 509026 434148
rect 509092 434136 509094 434148
rect 509094 434136 509126 434148
rect 508892 434114 508926 434136
rect 508992 434114 509026 434136
rect 509092 434114 509126 434136
rect 509192 434114 509226 434148
rect 509292 434114 509326 434148
rect 509392 434136 509420 434148
rect 509420 434136 509426 434148
rect 509392 434114 509426 434136
rect 508892 434046 508914 434048
rect 508914 434046 508926 434048
rect 508992 434046 509004 434048
rect 509004 434046 509026 434048
rect 509092 434046 509094 434048
rect 509094 434046 509126 434048
rect 508892 434014 508926 434046
rect 508992 434014 509026 434046
rect 509092 434014 509126 434046
rect 509192 434014 509226 434048
rect 509292 434014 509326 434048
rect 509392 434046 509420 434048
rect 509420 434046 509426 434048
rect 509392 434014 509426 434046
rect 508892 433914 508926 433948
rect 508992 433914 509026 433948
rect 509092 433914 509126 433948
rect 509192 433914 509226 433948
rect 509292 433914 509326 433948
rect 509392 433914 509426 433948
rect 508892 433814 508926 433848
rect 508992 433814 509026 433848
rect 509092 433814 509126 433848
rect 509192 433814 509226 433848
rect 509292 433814 509326 433848
rect 509392 433814 509426 433848
rect 508892 433720 508926 433748
rect 508992 433720 509026 433748
rect 509092 433720 509126 433748
rect 508892 433714 508914 433720
rect 508914 433714 508926 433720
rect 508992 433714 509004 433720
rect 509004 433714 509026 433720
rect 509092 433714 509094 433720
rect 509094 433714 509126 433720
rect 509192 433714 509226 433748
rect 509292 433714 509326 433748
rect 509392 433720 509426 433748
rect 509392 433714 509420 433720
rect 509420 433714 509426 433720
rect 510180 434226 510202 434248
rect 510202 434226 510214 434248
rect 510280 434226 510292 434248
rect 510292 434226 510314 434248
rect 510380 434226 510382 434248
rect 510382 434226 510414 434248
rect 510180 434214 510214 434226
rect 510280 434214 510314 434226
rect 510380 434214 510414 434226
rect 510480 434214 510514 434248
rect 510580 434214 510614 434248
rect 510680 434226 510708 434248
rect 510708 434226 510714 434248
rect 510680 434214 510714 434226
rect 510180 434136 510202 434148
rect 510202 434136 510214 434148
rect 510280 434136 510292 434148
rect 510292 434136 510314 434148
rect 510380 434136 510382 434148
rect 510382 434136 510414 434148
rect 510180 434114 510214 434136
rect 510280 434114 510314 434136
rect 510380 434114 510414 434136
rect 510480 434114 510514 434148
rect 510580 434114 510614 434148
rect 510680 434136 510708 434148
rect 510708 434136 510714 434148
rect 510680 434114 510714 434136
rect 510180 434046 510202 434048
rect 510202 434046 510214 434048
rect 510280 434046 510292 434048
rect 510292 434046 510314 434048
rect 510380 434046 510382 434048
rect 510382 434046 510414 434048
rect 510180 434014 510214 434046
rect 510280 434014 510314 434046
rect 510380 434014 510414 434046
rect 510480 434014 510514 434048
rect 510580 434014 510614 434048
rect 510680 434046 510708 434048
rect 510708 434046 510714 434048
rect 510680 434014 510714 434046
rect 510180 433914 510214 433948
rect 510280 433914 510314 433948
rect 510380 433914 510414 433948
rect 510480 433914 510514 433948
rect 510580 433914 510614 433948
rect 510680 433914 510714 433948
rect 510180 433814 510214 433848
rect 510280 433814 510314 433848
rect 510380 433814 510414 433848
rect 510480 433814 510514 433848
rect 510580 433814 510614 433848
rect 510680 433814 510714 433848
rect 510180 433720 510214 433748
rect 510280 433720 510314 433748
rect 510380 433720 510414 433748
rect 510180 433714 510202 433720
rect 510202 433714 510214 433720
rect 510280 433714 510292 433720
rect 510292 433714 510314 433720
rect 510380 433714 510382 433720
rect 510382 433714 510414 433720
rect 510480 433714 510514 433748
rect 510580 433714 510614 433748
rect 510680 433720 510714 433748
rect 510680 433714 510708 433720
rect 510708 433714 510714 433720
rect 511468 434226 511490 434248
rect 511490 434226 511502 434248
rect 511568 434226 511580 434248
rect 511580 434226 511602 434248
rect 511668 434226 511670 434248
rect 511670 434226 511702 434248
rect 511468 434214 511502 434226
rect 511568 434214 511602 434226
rect 511668 434214 511702 434226
rect 511768 434214 511802 434248
rect 511868 434214 511902 434248
rect 511968 434226 511996 434248
rect 511996 434226 512002 434248
rect 511968 434214 512002 434226
rect 511468 434136 511490 434148
rect 511490 434136 511502 434148
rect 511568 434136 511580 434148
rect 511580 434136 511602 434148
rect 511668 434136 511670 434148
rect 511670 434136 511702 434148
rect 511468 434114 511502 434136
rect 511568 434114 511602 434136
rect 511668 434114 511702 434136
rect 511768 434114 511802 434148
rect 511868 434114 511902 434148
rect 511968 434136 511996 434148
rect 511996 434136 512002 434148
rect 511968 434114 512002 434136
rect 511468 434046 511490 434048
rect 511490 434046 511502 434048
rect 511568 434046 511580 434048
rect 511580 434046 511602 434048
rect 511668 434046 511670 434048
rect 511670 434046 511702 434048
rect 511468 434014 511502 434046
rect 511568 434014 511602 434046
rect 511668 434014 511702 434046
rect 511768 434014 511802 434048
rect 511868 434014 511902 434048
rect 511968 434046 511996 434048
rect 511996 434046 512002 434048
rect 511968 434014 512002 434046
rect 511468 433914 511502 433948
rect 511568 433914 511602 433948
rect 511668 433914 511702 433948
rect 511768 433914 511802 433948
rect 511868 433914 511902 433948
rect 511968 433914 512002 433948
rect 511468 433814 511502 433848
rect 511568 433814 511602 433848
rect 511668 433814 511702 433848
rect 511768 433814 511802 433848
rect 511868 433814 511902 433848
rect 511968 433814 512002 433848
rect 511468 433720 511502 433748
rect 511568 433720 511602 433748
rect 511668 433720 511702 433748
rect 511468 433714 511490 433720
rect 511490 433714 511502 433720
rect 511568 433714 511580 433720
rect 511580 433714 511602 433720
rect 511668 433714 511670 433720
rect 511670 433714 511702 433720
rect 511768 433714 511802 433748
rect 511868 433714 511902 433748
rect 511968 433720 512002 433748
rect 511968 433714 511996 433720
rect 511996 433714 512002 433720
rect 512756 434226 512778 434248
rect 512778 434226 512790 434248
rect 512856 434226 512868 434248
rect 512868 434226 512890 434248
rect 512956 434226 512958 434248
rect 512958 434226 512990 434248
rect 512756 434214 512790 434226
rect 512856 434214 512890 434226
rect 512956 434214 512990 434226
rect 513056 434214 513090 434248
rect 513156 434214 513190 434248
rect 513256 434226 513284 434248
rect 513284 434226 513290 434248
rect 513256 434214 513290 434226
rect 512756 434136 512778 434148
rect 512778 434136 512790 434148
rect 512856 434136 512868 434148
rect 512868 434136 512890 434148
rect 512956 434136 512958 434148
rect 512958 434136 512990 434148
rect 512756 434114 512790 434136
rect 512856 434114 512890 434136
rect 512956 434114 512990 434136
rect 513056 434114 513090 434148
rect 513156 434114 513190 434148
rect 513256 434136 513284 434148
rect 513284 434136 513290 434148
rect 513256 434114 513290 434136
rect 512756 434046 512778 434048
rect 512778 434046 512790 434048
rect 512856 434046 512868 434048
rect 512868 434046 512890 434048
rect 512956 434046 512958 434048
rect 512958 434046 512990 434048
rect 512756 434014 512790 434046
rect 512856 434014 512890 434046
rect 512956 434014 512990 434046
rect 513056 434014 513090 434048
rect 513156 434014 513190 434048
rect 513256 434046 513284 434048
rect 513284 434046 513290 434048
rect 513256 434014 513290 434046
rect 512756 433914 512790 433948
rect 512856 433914 512890 433948
rect 512956 433914 512990 433948
rect 513056 433914 513090 433948
rect 513156 433914 513190 433948
rect 513256 433914 513290 433948
rect 512756 433814 512790 433848
rect 512856 433814 512890 433848
rect 512956 433814 512990 433848
rect 513056 433814 513090 433848
rect 513156 433814 513190 433848
rect 513256 433814 513290 433848
rect 512756 433720 512790 433748
rect 512856 433720 512890 433748
rect 512956 433720 512990 433748
rect 512756 433714 512778 433720
rect 512778 433714 512790 433720
rect 512856 433714 512868 433720
rect 512868 433714 512890 433720
rect 512956 433714 512958 433720
rect 512958 433714 512990 433720
rect 513056 433714 513090 433748
rect 513156 433714 513190 433748
rect 513256 433720 513290 433748
rect 513256 433714 513284 433720
rect 513284 433714 513290 433720
rect 500418 433408 500518 433508
rect 500642 433408 500742 433508
rect 500866 433408 500966 433508
rect 501090 433408 501190 433508
rect 501314 433408 501368 433508
rect 501368 433408 501414 433508
rect 500418 433184 500518 433284
rect 500642 433184 500742 433284
rect 500866 433184 500966 433284
rect 501090 433184 501190 433284
rect 501314 433184 501368 433284
rect 501368 433184 501414 433284
rect 500418 432960 500518 433060
rect 500642 432960 500742 433060
rect 500866 432960 500966 433060
rect 501090 432960 501190 433060
rect 501314 432960 501368 433060
rect 501368 432960 501414 433060
rect 500418 432736 500518 432836
rect 500642 432736 500742 432836
rect 500866 432736 500966 432836
rect 501090 432736 501190 432836
rect 501314 432736 501368 432836
rect 501368 432736 501414 432836
rect 500418 432512 500518 432612
rect 500642 432512 500742 432612
rect 500866 432512 500966 432612
rect 501090 432512 501190 432612
rect 501314 432512 501368 432612
rect 501368 432512 501414 432612
rect 500418 432288 500518 432388
rect 500642 432288 500742 432388
rect 500866 432288 500966 432388
rect 501090 432288 501190 432388
rect 501314 432288 501368 432388
rect 501368 432288 501414 432388
rect 503740 432938 503762 432960
rect 503762 432938 503774 432960
rect 503840 432938 503852 432960
rect 503852 432938 503874 432960
rect 503940 432938 503942 432960
rect 503942 432938 503974 432960
rect 503740 432926 503774 432938
rect 503840 432926 503874 432938
rect 503940 432926 503974 432938
rect 504040 432926 504074 432960
rect 504140 432926 504174 432960
rect 504240 432938 504268 432960
rect 504268 432938 504274 432960
rect 504240 432926 504274 432938
rect 503740 432848 503762 432860
rect 503762 432848 503774 432860
rect 503840 432848 503852 432860
rect 503852 432848 503874 432860
rect 503940 432848 503942 432860
rect 503942 432848 503974 432860
rect 503740 432826 503774 432848
rect 503840 432826 503874 432848
rect 503940 432826 503974 432848
rect 504040 432826 504074 432860
rect 504140 432826 504174 432860
rect 504240 432848 504268 432860
rect 504268 432848 504274 432860
rect 504240 432826 504274 432848
rect 503740 432758 503762 432760
rect 503762 432758 503774 432760
rect 503840 432758 503852 432760
rect 503852 432758 503874 432760
rect 503940 432758 503942 432760
rect 503942 432758 503974 432760
rect 503740 432726 503774 432758
rect 503840 432726 503874 432758
rect 503940 432726 503974 432758
rect 504040 432726 504074 432760
rect 504140 432726 504174 432760
rect 504240 432758 504268 432760
rect 504268 432758 504274 432760
rect 504240 432726 504274 432758
rect 503740 432626 503774 432660
rect 503840 432626 503874 432660
rect 503940 432626 503974 432660
rect 504040 432626 504074 432660
rect 504140 432626 504174 432660
rect 504240 432626 504274 432660
rect 503740 432526 503774 432560
rect 503840 432526 503874 432560
rect 503940 432526 503974 432560
rect 504040 432526 504074 432560
rect 504140 432526 504174 432560
rect 504240 432526 504274 432560
rect 503740 432432 503774 432460
rect 503840 432432 503874 432460
rect 503940 432432 503974 432460
rect 503740 432426 503762 432432
rect 503762 432426 503774 432432
rect 503840 432426 503852 432432
rect 503852 432426 503874 432432
rect 503940 432426 503942 432432
rect 503942 432426 503974 432432
rect 504040 432426 504074 432460
rect 504140 432426 504174 432460
rect 504240 432432 504274 432460
rect 504240 432426 504268 432432
rect 504268 432426 504274 432432
rect 505028 432938 505050 432960
rect 505050 432938 505062 432960
rect 505128 432938 505140 432960
rect 505140 432938 505162 432960
rect 505228 432938 505230 432960
rect 505230 432938 505262 432960
rect 505028 432926 505062 432938
rect 505128 432926 505162 432938
rect 505228 432926 505262 432938
rect 505328 432926 505362 432960
rect 505428 432926 505462 432960
rect 505528 432938 505556 432960
rect 505556 432938 505562 432960
rect 505528 432926 505562 432938
rect 505028 432848 505050 432860
rect 505050 432848 505062 432860
rect 505128 432848 505140 432860
rect 505140 432848 505162 432860
rect 505228 432848 505230 432860
rect 505230 432848 505262 432860
rect 505028 432826 505062 432848
rect 505128 432826 505162 432848
rect 505228 432826 505262 432848
rect 505328 432826 505362 432860
rect 505428 432826 505462 432860
rect 505528 432848 505556 432860
rect 505556 432848 505562 432860
rect 505528 432826 505562 432848
rect 505028 432758 505050 432760
rect 505050 432758 505062 432760
rect 505128 432758 505140 432760
rect 505140 432758 505162 432760
rect 505228 432758 505230 432760
rect 505230 432758 505262 432760
rect 505028 432726 505062 432758
rect 505128 432726 505162 432758
rect 505228 432726 505262 432758
rect 505328 432726 505362 432760
rect 505428 432726 505462 432760
rect 505528 432758 505556 432760
rect 505556 432758 505562 432760
rect 505528 432726 505562 432758
rect 505028 432626 505062 432660
rect 505128 432626 505162 432660
rect 505228 432626 505262 432660
rect 505328 432626 505362 432660
rect 505428 432626 505462 432660
rect 505528 432626 505562 432660
rect 505028 432526 505062 432560
rect 505128 432526 505162 432560
rect 505228 432526 505262 432560
rect 505328 432526 505362 432560
rect 505428 432526 505462 432560
rect 505528 432526 505562 432560
rect 505028 432432 505062 432460
rect 505128 432432 505162 432460
rect 505228 432432 505262 432460
rect 505028 432426 505050 432432
rect 505050 432426 505062 432432
rect 505128 432426 505140 432432
rect 505140 432426 505162 432432
rect 505228 432426 505230 432432
rect 505230 432426 505262 432432
rect 505328 432426 505362 432460
rect 505428 432426 505462 432460
rect 505528 432432 505562 432460
rect 505528 432426 505556 432432
rect 505556 432426 505562 432432
rect 506316 432938 506338 432960
rect 506338 432938 506350 432960
rect 506416 432938 506428 432960
rect 506428 432938 506450 432960
rect 506516 432938 506518 432960
rect 506518 432938 506550 432960
rect 506316 432926 506350 432938
rect 506416 432926 506450 432938
rect 506516 432926 506550 432938
rect 506616 432926 506650 432960
rect 506716 432926 506750 432960
rect 506816 432938 506844 432960
rect 506844 432938 506850 432960
rect 506816 432926 506850 432938
rect 506316 432848 506338 432860
rect 506338 432848 506350 432860
rect 506416 432848 506428 432860
rect 506428 432848 506450 432860
rect 506516 432848 506518 432860
rect 506518 432848 506550 432860
rect 506316 432826 506350 432848
rect 506416 432826 506450 432848
rect 506516 432826 506550 432848
rect 506616 432826 506650 432860
rect 506716 432826 506750 432860
rect 506816 432848 506844 432860
rect 506844 432848 506850 432860
rect 506816 432826 506850 432848
rect 506316 432758 506338 432760
rect 506338 432758 506350 432760
rect 506416 432758 506428 432760
rect 506428 432758 506450 432760
rect 506516 432758 506518 432760
rect 506518 432758 506550 432760
rect 506316 432726 506350 432758
rect 506416 432726 506450 432758
rect 506516 432726 506550 432758
rect 506616 432726 506650 432760
rect 506716 432726 506750 432760
rect 506816 432758 506844 432760
rect 506844 432758 506850 432760
rect 506816 432726 506850 432758
rect 506316 432626 506350 432660
rect 506416 432626 506450 432660
rect 506516 432626 506550 432660
rect 506616 432626 506650 432660
rect 506716 432626 506750 432660
rect 506816 432626 506850 432660
rect 506316 432526 506350 432560
rect 506416 432526 506450 432560
rect 506516 432526 506550 432560
rect 506616 432526 506650 432560
rect 506716 432526 506750 432560
rect 506816 432526 506850 432560
rect 506316 432432 506350 432460
rect 506416 432432 506450 432460
rect 506516 432432 506550 432460
rect 506316 432426 506338 432432
rect 506338 432426 506350 432432
rect 506416 432426 506428 432432
rect 506428 432426 506450 432432
rect 506516 432426 506518 432432
rect 506518 432426 506550 432432
rect 506616 432426 506650 432460
rect 506716 432426 506750 432460
rect 506816 432432 506850 432460
rect 506816 432426 506844 432432
rect 506844 432426 506850 432432
rect 507604 432938 507626 432960
rect 507626 432938 507638 432960
rect 507704 432938 507716 432960
rect 507716 432938 507738 432960
rect 507804 432938 507806 432960
rect 507806 432938 507838 432960
rect 507604 432926 507638 432938
rect 507704 432926 507738 432938
rect 507804 432926 507838 432938
rect 507904 432926 507938 432960
rect 508004 432926 508038 432960
rect 508104 432938 508132 432960
rect 508132 432938 508138 432960
rect 508104 432926 508138 432938
rect 507604 432848 507626 432860
rect 507626 432848 507638 432860
rect 507704 432848 507716 432860
rect 507716 432848 507738 432860
rect 507804 432848 507806 432860
rect 507806 432848 507838 432860
rect 507604 432826 507638 432848
rect 507704 432826 507738 432848
rect 507804 432826 507838 432848
rect 507904 432826 507938 432860
rect 508004 432826 508038 432860
rect 508104 432848 508132 432860
rect 508132 432848 508138 432860
rect 508104 432826 508138 432848
rect 507604 432758 507626 432760
rect 507626 432758 507638 432760
rect 507704 432758 507716 432760
rect 507716 432758 507738 432760
rect 507804 432758 507806 432760
rect 507806 432758 507838 432760
rect 507604 432726 507638 432758
rect 507704 432726 507738 432758
rect 507804 432726 507838 432758
rect 507904 432726 507938 432760
rect 508004 432726 508038 432760
rect 508104 432758 508132 432760
rect 508132 432758 508138 432760
rect 508104 432726 508138 432758
rect 507604 432626 507638 432660
rect 507704 432626 507738 432660
rect 507804 432626 507838 432660
rect 507904 432626 507938 432660
rect 508004 432626 508038 432660
rect 508104 432626 508138 432660
rect 507604 432526 507638 432560
rect 507704 432526 507738 432560
rect 507804 432526 507838 432560
rect 507904 432526 507938 432560
rect 508004 432526 508038 432560
rect 508104 432526 508138 432560
rect 507604 432432 507638 432460
rect 507704 432432 507738 432460
rect 507804 432432 507838 432460
rect 507604 432426 507626 432432
rect 507626 432426 507638 432432
rect 507704 432426 507716 432432
rect 507716 432426 507738 432432
rect 507804 432426 507806 432432
rect 507806 432426 507838 432432
rect 507904 432426 507938 432460
rect 508004 432426 508038 432460
rect 508104 432432 508138 432460
rect 508104 432426 508132 432432
rect 508132 432426 508138 432432
rect 508892 432938 508914 432960
rect 508914 432938 508926 432960
rect 508992 432938 509004 432960
rect 509004 432938 509026 432960
rect 509092 432938 509094 432960
rect 509094 432938 509126 432960
rect 508892 432926 508926 432938
rect 508992 432926 509026 432938
rect 509092 432926 509126 432938
rect 509192 432926 509226 432960
rect 509292 432926 509326 432960
rect 509392 432938 509420 432960
rect 509420 432938 509426 432960
rect 509392 432926 509426 432938
rect 508892 432848 508914 432860
rect 508914 432848 508926 432860
rect 508992 432848 509004 432860
rect 509004 432848 509026 432860
rect 509092 432848 509094 432860
rect 509094 432848 509126 432860
rect 508892 432826 508926 432848
rect 508992 432826 509026 432848
rect 509092 432826 509126 432848
rect 509192 432826 509226 432860
rect 509292 432826 509326 432860
rect 509392 432848 509420 432860
rect 509420 432848 509426 432860
rect 509392 432826 509426 432848
rect 508892 432758 508914 432760
rect 508914 432758 508926 432760
rect 508992 432758 509004 432760
rect 509004 432758 509026 432760
rect 509092 432758 509094 432760
rect 509094 432758 509126 432760
rect 508892 432726 508926 432758
rect 508992 432726 509026 432758
rect 509092 432726 509126 432758
rect 509192 432726 509226 432760
rect 509292 432726 509326 432760
rect 509392 432758 509420 432760
rect 509420 432758 509426 432760
rect 509392 432726 509426 432758
rect 508892 432626 508926 432660
rect 508992 432626 509026 432660
rect 509092 432626 509126 432660
rect 509192 432626 509226 432660
rect 509292 432626 509326 432660
rect 509392 432626 509426 432660
rect 508892 432526 508926 432560
rect 508992 432526 509026 432560
rect 509092 432526 509126 432560
rect 509192 432526 509226 432560
rect 509292 432526 509326 432560
rect 509392 432526 509426 432560
rect 508892 432432 508926 432460
rect 508992 432432 509026 432460
rect 509092 432432 509126 432460
rect 508892 432426 508914 432432
rect 508914 432426 508926 432432
rect 508992 432426 509004 432432
rect 509004 432426 509026 432432
rect 509092 432426 509094 432432
rect 509094 432426 509126 432432
rect 509192 432426 509226 432460
rect 509292 432426 509326 432460
rect 509392 432432 509426 432460
rect 509392 432426 509420 432432
rect 509420 432426 509426 432432
rect 510180 432938 510202 432960
rect 510202 432938 510214 432960
rect 510280 432938 510292 432960
rect 510292 432938 510314 432960
rect 510380 432938 510382 432960
rect 510382 432938 510414 432960
rect 510180 432926 510214 432938
rect 510280 432926 510314 432938
rect 510380 432926 510414 432938
rect 510480 432926 510514 432960
rect 510580 432926 510614 432960
rect 510680 432938 510708 432960
rect 510708 432938 510714 432960
rect 510680 432926 510714 432938
rect 510180 432848 510202 432860
rect 510202 432848 510214 432860
rect 510280 432848 510292 432860
rect 510292 432848 510314 432860
rect 510380 432848 510382 432860
rect 510382 432848 510414 432860
rect 510180 432826 510214 432848
rect 510280 432826 510314 432848
rect 510380 432826 510414 432848
rect 510480 432826 510514 432860
rect 510580 432826 510614 432860
rect 510680 432848 510708 432860
rect 510708 432848 510714 432860
rect 510680 432826 510714 432848
rect 510180 432758 510202 432760
rect 510202 432758 510214 432760
rect 510280 432758 510292 432760
rect 510292 432758 510314 432760
rect 510380 432758 510382 432760
rect 510382 432758 510414 432760
rect 510180 432726 510214 432758
rect 510280 432726 510314 432758
rect 510380 432726 510414 432758
rect 510480 432726 510514 432760
rect 510580 432726 510614 432760
rect 510680 432758 510708 432760
rect 510708 432758 510714 432760
rect 510680 432726 510714 432758
rect 510180 432626 510214 432660
rect 510280 432626 510314 432660
rect 510380 432626 510414 432660
rect 510480 432626 510514 432660
rect 510580 432626 510614 432660
rect 510680 432626 510714 432660
rect 510180 432526 510214 432560
rect 510280 432526 510314 432560
rect 510380 432526 510414 432560
rect 510480 432526 510514 432560
rect 510580 432526 510614 432560
rect 510680 432526 510714 432560
rect 510180 432432 510214 432460
rect 510280 432432 510314 432460
rect 510380 432432 510414 432460
rect 510180 432426 510202 432432
rect 510202 432426 510214 432432
rect 510280 432426 510292 432432
rect 510292 432426 510314 432432
rect 510380 432426 510382 432432
rect 510382 432426 510414 432432
rect 510480 432426 510514 432460
rect 510580 432426 510614 432460
rect 510680 432432 510714 432460
rect 510680 432426 510708 432432
rect 510708 432426 510714 432432
rect 511468 432938 511490 432960
rect 511490 432938 511502 432960
rect 511568 432938 511580 432960
rect 511580 432938 511602 432960
rect 511668 432938 511670 432960
rect 511670 432938 511702 432960
rect 511468 432926 511502 432938
rect 511568 432926 511602 432938
rect 511668 432926 511702 432938
rect 511768 432926 511802 432960
rect 511868 432926 511902 432960
rect 511968 432938 511996 432960
rect 511996 432938 512002 432960
rect 511968 432926 512002 432938
rect 511468 432848 511490 432860
rect 511490 432848 511502 432860
rect 511568 432848 511580 432860
rect 511580 432848 511602 432860
rect 511668 432848 511670 432860
rect 511670 432848 511702 432860
rect 511468 432826 511502 432848
rect 511568 432826 511602 432848
rect 511668 432826 511702 432848
rect 511768 432826 511802 432860
rect 511868 432826 511902 432860
rect 511968 432848 511996 432860
rect 511996 432848 512002 432860
rect 511968 432826 512002 432848
rect 511468 432758 511490 432760
rect 511490 432758 511502 432760
rect 511568 432758 511580 432760
rect 511580 432758 511602 432760
rect 511668 432758 511670 432760
rect 511670 432758 511702 432760
rect 511468 432726 511502 432758
rect 511568 432726 511602 432758
rect 511668 432726 511702 432758
rect 511768 432726 511802 432760
rect 511868 432726 511902 432760
rect 511968 432758 511996 432760
rect 511996 432758 512002 432760
rect 511968 432726 512002 432758
rect 511468 432626 511502 432660
rect 511568 432626 511602 432660
rect 511668 432626 511702 432660
rect 511768 432626 511802 432660
rect 511868 432626 511902 432660
rect 511968 432626 512002 432660
rect 511468 432526 511502 432560
rect 511568 432526 511602 432560
rect 511668 432526 511702 432560
rect 511768 432526 511802 432560
rect 511868 432526 511902 432560
rect 511968 432526 512002 432560
rect 511468 432432 511502 432460
rect 511568 432432 511602 432460
rect 511668 432432 511702 432460
rect 511468 432426 511490 432432
rect 511490 432426 511502 432432
rect 511568 432426 511580 432432
rect 511580 432426 511602 432432
rect 511668 432426 511670 432432
rect 511670 432426 511702 432432
rect 511768 432426 511802 432460
rect 511868 432426 511902 432460
rect 511968 432432 512002 432460
rect 511968 432426 511996 432432
rect 511996 432426 512002 432432
rect 512756 432938 512778 432960
rect 512778 432938 512790 432960
rect 512856 432938 512868 432960
rect 512868 432938 512890 432960
rect 512956 432938 512958 432960
rect 512958 432938 512990 432960
rect 512756 432926 512790 432938
rect 512856 432926 512890 432938
rect 512956 432926 512990 432938
rect 513056 432926 513090 432960
rect 513156 432926 513190 432960
rect 513256 432938 513284 432960
rect 513284 432938 513290 432960
rect 513256 432926 513290 432938
rect 512756 432848 512778 432860
rect 512778 432848 512790 432860
rect 512856 432848 512868 432860
rect 512868 432848 512890 432860
rect 512956 432848 512958 432860
rect 512958 432848 512990 432860
rect 512756 432826 512790 432848
rect 512856 432826 512890 432848
rect 512956 432826 512990 432848
rect 513056 432826 513090 432860
rect 513156 432826 513190 432860
rect 513256 432848 513284 432860
rect 513284 432848 513290 432860
rect 513256 432826 513290 432848
rect 512756 432758 512778 432760
rect 512778 432758 512790 432760
rect 512856 432758 512868 432760
rect 512868 432758 512890 432760
rect 512956 432758 512958 432760
rect 512958 432758 512990 432760
rect 512756 432726 512790 432758
rect 512856 432726 512890 432758
rect 512956 432726 512990 432758
rect 513056 432726 513090 432760
rect 513156 432726 513190 432760
rect 513256 432758 513284 432760
rect 513284 432758 513290 432760
rect 513256 432726 513290 432758
rect 512756 432626 512790 432660
rect 512856 432626 512890 432660
rect 512956 432626 512990 432660
rect 513056 432626 513090 432660
rect 513156 432626 513190 432660
rect 513256 432626 513290 432660
rect 512756 432526 512790 432560
rect 512856 432526 512890 432560
rect 512956 432526 512990 432560
rect 513056 432526 513090 432560
rect 513156 432526 513190 432560
rect 513256 432526 513290 432560
rect 512756 432432 512790 432460
rect 512856 432432 512890 432460
rect 512956 432432 512990 432460
rect 512756 432426 512778 432432
rect 512778 432426 512790 432432
rect 512856 432426 512868 432432
rect 512868 432426 512890 432432
rect 512956 432426 512958 432432
rect 512958 432426 512990 432432
rect 513056 432426 513090 432460
rect 513156 432426 513190 432460
rect 513256 432432 513290 432460
rect 513256 432426 513284 432432
rect 513284 432426 513290 432432
rect 500418 432068 500518 432164
rect 500642 432068 500742 432164
rect 500866 432068 500966 432164
rect 501090 432068 501190 432164
rect 501314 432068 501368 432164
rect 501368 432068 501414 432164
rect 500418 432064 500518 432068
rect 500642 432064 500742 432068
rect 500866 432064 500966 432068
rect 501090 432064 501190 432068
rect 501314 432064 501414 432068
rect 500418 431840 500518 431940
rect 500642 431840 500742 431940
rect 500866 431840 500966 431940
rect 501090 431840 501190 431940
rect 501314 431840 501414 431940
rect 500418 431616 500518 431716
rect 500642 431616 500742 431716
rect 500866 431616 500966 431716
rect 501090 431616 501190 431716
rect 501314 431616 501414 431716
rect 500418 431392 500518 431492
rect 500642 431392 500742 431492
rect 500866 431392 500966 431492
rect 501090 431392 501190 431492
rect 501314 431392 501414 431492
rect 500418 431168 500518 431268
rect 500642 431168 500742 431268
rect 500866 431168 500966 431268
rect 501090 431168 501190 431268
rect 501314 431168 501414 431268
rect 500418 430944 500518 431044
rect 500642 430944 500742 431044
rect 500866 430944 500966 431044
rect 501090 430944 501190 431044
rect 501314 430944 501414 431044
rect 503920 430926 504020 431026
rect 504144 430926 504244 431026
rect 504368 430926 504468 431026
rect 504592 430926 504692 431026
rect 504816 430926 504916 431026
rect 505040 430926 505140 431026
rect 505264 430926 505364 431026
rect 505488 430926 505588 431026
rect 505712 430926 505812 431026
rect 505936 430926 506036 431026
rect 506160 430926 506260 431026
rect 506384 430926 506484 431026
rect 506608 430926 506708 431026
rect 506832 430926 506932 431026
rect 507056 430926 507156 431026
rect 507280 430926 507380 431026
rect 507504 430926 507604 431026
rect 507728 430926 507828 431026
rect 507952 430926 508052 431026
rect 508176 430926 508276 431026
rect 508400 430926 508500 431026
rect 508624 430926 508724 431026
rect 508848 430926 508948 431026
rect 509072 430926 509172 431026
rect 509296 430926 509396 431026
rect 509520 430926 509620 431026
rect 509744 430926 509844 431026
rect 509968 430926 510068 431026
rect 510192 430926 510292 431026
rect 510416 430926 510516 431026
rect 517320 430926 517420 431026
rect 517544 430926 517644 431026
rect 517768 430926 517868 431026
rect 517992 430926 518092 431026
rect 518216 430926 518316 431026
rect 518440 430926 518540 431026
rect 518664 430926 518764 431026
rect 518888 430926 518988 431026
rect 519112 430926 519212 431026
rect 519336 430926 519436 431026
rect 519560 430926 519660 431026
rect 519784 430926 519884 431026
rect 520008 430926 520108 431026
rect 520232 430926 520332 431026
rect 520456 430926 520556 431026
rect 520680 430926 520780 431026
rect 520904 430926 521004 431026
rect 521128 430926 521228 431026
rect 521352 430926 521452 431026
rect 521576 430926 521676 431026
rect 521800 430926 521900 431026
rect 522024 430926 522124 431026
rect 522248 430926 522348 431026
rect 522472 430926 522572 431026
rect 522696 430926 522796 431026
rect 522920 430926 523020 431026
rect 523144 430926 523244 431026
rect 523368 430926 523468 431026
rect 523592 430926 523692 431026
rect 523816 430926 523916 431026
rect 527618 474180 527718 474280
rect 527842 474180 527942 474280
rect 528066 474180 528166 474280
rect 528290 474180 528390 474280
rect 528514 474180 528592 474280
rect 528592 474180 528614 474280
rect 527618 473956 527718 474056
rect 527842 473956 527942 474056
rect 528066 473956 528166 474056
rect 528290 473956 528390 474056
rect 528514 473956 528592 474056
rect 528592 473956 528614 474056
rect 527618 473732 527718 473832
rect 527842 473732 527942 473832
rect 528066 473732 528166 473832
rect 528290 473732 528390 473832
rect 528514 473732 528592 473832
rect 528592 473732 528614 473832
rect 527618 473508 527718 473608
rect 527842 473508 527942 473608
rect 528066 473508 528166 473608
rect 528290 473508 528390 473608
rect 528514 473508 528592 473608
rect 528592 473508 528614 473608
rect 527618 473284 527718 473384
rect 527842 473284 527942 473384
rect 528066 473284 528166 473384
rect 528290 473284 528390 473384
rect 528514 473284 528592 473384
rect 528592 473284 528614 473384
rect 527618 473060 527718 473160
rect 527842 473060 527942 473160
rect 528066 473060 528166 473160
rect 528290 473060 528390 473160
rect 528514 473060 528592 473160
rect 528592 473060 528614 473160
rect 527618 472836 527718 472936
rect 527842 472836 527942 472936
rect 528066 472836 528166 472936
rect 528290 472836 528390 472936
rect 528514 472836 528592 472936
rect 528592 472836 528614 472936
rect 527618 472612 527718 472712
rect 527842 472612 527942 472712
rect 528066 472612 528166 472712
rect 528290 472612 528390 472712
rect 528514 472612 528592 472712
rect 528592 472612 528614 472712
rect 527618 472388 527718 472488
rect 527842 472388 527942 472488
rect 528066 472388 528166 472488
rect 528290 472388 528390 472488
rect 528514 472388 528592 472488
rect 528592 472388 528614 472488
rect 527618 472164 527718 472264
rect 527842 472164 527942 472264
rect 528066 472164 528166 472264
rect 528290 472164 528390 472264
rect 528514 472164 528592 472264
rect 528592 472164 528614 472264
rect 527618 471940 527718 472040
rect 527842 471940 527942 472040
rect 528066 471940 528166 472040
rect 528290 471940 528390 472040
rect 528514 471940 528592 472040
rect 528592 471940 528614 472040
rect 527618 471716 527718 471816
rect 527842 471716 527942 471816
rect 528066 471716 528166 471816
rect 528290 471716 528390 471816
rect 528514 471716 528592 471816
rect 528592 471716 528614 471816
rect 527618 471492 527718 471592
rect 527842 471492 527942 471592
rect 528066 471492 528166 471592
rect 528290 471492 528390 471592
rect 528514 471492 528592 471592
rect 528592 471492 528614 471592
rect 527618 471268 527718 471368
rect 527842 471268 527942 471368
rect 528066 471268 528166 471368
rect 528290 471268 528390 471368
rect 528514 471268 528592 471368
rect 528592 471268 528614 471368
rect 527618 471044 527718 471144
rect 527842 471044 527942 471144
rect 528066 471044 528166 471144
rect 528290 471044 528390 471144
rect 528514 471044 528592 471144
rect 528592 471044 528614 471144
rect 527618 470820 527718 470920
rect 527842 470820 527942 470920
rect 528066 470820 528166 470920
rect 528290 470820 528390 470920
rect 528514 470820 528592 470920
rect 528592 470820 528614 470920
rect 527618 470596 527718 470696
rect 527842 470596 527942 470696
rect 528066 470596 528166 470696
rect 528290 470596 528390 470696
rect 528514 470596 528592 470696
rect 528592 470596 528614 470696
rect 527618 470372 527718 470472
rect 527842 470372 527942 470472
rect 528066 470372 528166 470472
rect 528290 470372 528390 470472
rect 528514 470372 528592 470472
rect 528592 470372 528614 470472
rect 527618 470148 527718 470248
rect 527842 470148 527942 470248
rect 528066 470148 528166 470248
rect 528290 470148 528390 470248
rect 528514 470148 528592 470248
rect 528592 470148 528614 470248
rect 527618 469924 527718 470024
rect 527842 469924 527942 470024
rect 528066 469924 528166 470024
rect 528290 469924 528390 470024
rect 528514 469924 528592 470024
rect 528592 469924 528614 470024
rect 527618 469700 527718 469800
rect 527842 469700 527942 469800
rect 528066 469700 528166 469800
rect 528290 469700 528390 469800
rect 528514 469700 528592 469800
rect 528592 469700 528614 469800
rect 527618 469476 527718 469576
rect 527842 469476 527942 469576
rect 528066 469476 528166 469576
rect 528290 469476 528390 469576
rect 528514 469476 528592 469576
rect 528592 469476 528614 469576
rect 527618 469252 527718 469352
rect 527842 469252 527942 469352
rect 528066 469252 528166 469352
rect 528290 469252 528390 469352
rect 528514 469252 528592 469352
rect 528592 469252 528614 469352
rect 527618 469028 527718 469128
rect 527842 469028 527942 469128
rect 528066 469028 528166 469128
rect 528290 469028 528390 469128
rect 528514 469028 528592 469128
rect 528592 469028 528614 469128
rect 527618 468804 527718 468904
rect 527842 468804 527942 468904
rect 528066 468804 528166 468904
rect 528290 468804 528390 468904
rect 528514 468804 528592 468904
rect 528592 468804 528614 468904
rect 527618 468580 527718 468680
rect 527842 468580 527942 468680
rect 528066 468580 528166 468680
rect 528290 468580 528390 468680
rect 528514 468580 528592 468680
rect 528592 468580 528614 468680
rect 527618 468356 527718 468456
rect 527842 468356 527942 468456
rect 528066 468356 528166 468456
rect 528290 468356 528390 468456
rect 528514 468356 528592 468456
rect 528592 468356 528614 468456
rect 527618 468132 527718 468232
rect 527842 468132 527942 468232
rect 528066 468132 528166 468232
rect 528290 468132 528390 468232
rect 528514 468132 528592 468232
rect 528592 468132 528614 468232
rect 527618 467908 527718 468008
rect 527842 467908 527942 468008
rect 528066 467908 528166 468008
rect 528290 467908 528390 468008
rect 528514 467908 528592 468008
rect 528592 467908 528614 468008
rect 527618 467684 527718 467784
rect 527842 467684 527942 467784
rect 528066 467684 528166 467784
rect 528290 467684 528390 467784
rect 528514 467684 528592 467784
rect 528592 467684 528614 467784
rect 527618 463710 527718 463810
rect 527842 463710 527942 463810
rect 528066 463710 528166 463810
rect 528290 463710 528390 463810
rect 528514 463710 528592 463810
rect 528592 463710 528614 463810
rect 527618 463486 527718 463586
rect 527842 463486 527942 463586
rect 528066 463486 528166 463586
rect 528290 463486 528390 463586
rect 528514 463486 528592 463586
rect 528592 463486 528614 463586
rect 527618 463262 527718 463362
rect 527842 463262 527942 463362
rect 528066 463262 528166 463362
rect 528290 463262 528390 463362
rect 528514 463262 528592 463362
rect 528592 463262 528614 463362
rect 527618 463038 527718 463138
rect 527842 463038 527942 463138
rect 528066 463038 528166 463138
rect 528290 463038 528390 463138
rect 528514 463038 528592 463138
rect 528592 463038 528614 463138
rect 527618 462814 527718 462914
rect 527842 462814 527942 462914
rect 528066 462814 528166 462914
rect 528290 462814 528390 462914
rect 528514 462814 528592 462914
rect 528592 462814 528614 462914
rect 527618 462590 527718 462690
rect 527842 462590 527942 462690
rect 528066 462590 528166 462690
rect 528290 462590 528390 462690
rect 528514 462590 528592 462690
rect 528592 462590 528614 462690
rect 527618 462366 527718 462466
rect 527842 462366 527942 462466
rect 528066 462366 528166 462466
rect 528290 462366 528390 462466
rect 528514 462366 528592 462466
rect 528592 462366 528614 462466
rect 527618 462142 527718 462242
rect 527842 462142 527942 462242
rect 528066 462142 528166 462242
rect 528290 462142 528390 462242
rect 528514 462142 528592 462242
rect 528592 462142 528614 462242
rect 527618 461918 527718 462018
rect 527842 461918 527942 462018
rect 528066 461918 528166 462018
rect 528290 461918 528390 462018
rect 528514 461918 528592 462018
rect 528592 461918 528614 462018
rect 527618 461694 527718 461794
rect 527842 461694 527942 461794
rect 528066 461694 528166 461794
rect 528290 461694 528390 461794
rect 528514 461694 528592 461794
rect 528592 461694 528614 461794
rect 527618 461470 527718 461570
rect 527842 461470 527942 461570
rect 528066 461470 528166 461570
rect 528290 461470 528390 461570
rect 528514 461470 528592 461570
rect 528592 461470 528614 461570
rect 527618 461246 527718 461346
rect 527842 461246 527942 461346
rect 528066 461246 528166 461346
rect 528290 461246 528390 461346
rect 528514 461246 528592 461346
rect 528592 461246 528614 461346
rect 527618 461022 527718 461122
rect 527842 461022 527942 461122
rect 528066 461022 528166 461122
rect 528290 461022 528390 461122
rect 528514 461022 528592 461122
rect 528592 461022 528614 461122
rect 527618 460798 527718 460898
rect 527842 460798 527942 460898
rect 528066 460798 528166 460898
rect 528290 460798 528390 460898
rect 528514 460798 528592 460898
rect 528592 460798 528614 460898
rect 527618 460574 527718 460674
rect 527842 460574 527942 460674
rect 528066 460574 528166 460674
rect 528290 460574 528390 460674
rect 528514 460574 528592 460674
rect 528592 460574 528614 460674
rect 527618 460350 527718 460450
rect 527842 460350 527942 460450
rect 528066 460350 528166 460450
rect 528290 460350 528390 460450
rect 528514 460350 528592 460450
rect 528592 460350 528614 460450
rect 527618 460126 527718 460226
rect 527842 460126 527942 460226
rect 528066 460126 528166 460226
rect 528290 460126 528390 460226
rect 528514 460126 528592 460226
rect 528592 460126 528614 460226
rect 527618 459902 527718 460002
rect 527842 459902 527942 460002
rect 528066 459902 528166 460002
rect 528290 459902 528390 460002
rect 528514 459902 528592 460002
rect 528592 459902 528614 460002
rect 527618 459678 527718 459778
rect 527842 459678 527942 459778
rect 528066 459678 528166 459778
rect 528290 459678 528390 459778
rect 528514 459678 528592 459778
rect 528592 459678 528614 459778
rect 527618 459454 527718 459554
rect 527842 459454 527942 459554
rect 528066 459454 528166 459554
rect 528290 459454 528390 459554
rect 528514 459454 528592 459554
rect 528592 459454 528614 459554
rect 527618 459230 527718 459330
rect 527842 459230 527942 459330
rect 528066 459230 528166 459330
rect 528290 459230 528390 459330
rect 528514 459230 528592 459330
rect 528592 459230 528614 459330
rect 527618 459006 527718 459106
rect 527842 459006 527942 459106
rect 528066 459006 528166 459106
rect 528290 459006 528390 459106
rect 528514 459006 528592 459106
rect 528592 459006 528614 459106
rect 527618 458782 527718 458882
rect 527842 458782 527942 458882
rect 528066 458782 528166 458882
rect 528290 458782 528390 458882
rect 528514 458782 528592 458882
rect 528592 458782 528614 458882
rect 527618 458558 527718 458658
rect 527842 458558 527942 458658
rect 528066 458558 528166 458658
rect 528290 458558 528390 458658
rect 528514 458558 528592 458658
rect 528592 458558 528614 458658
rect 527618 458334 527718 458434
rect 527842 458334 527942 458434
rect 528066 458334 528166 458434
rect 528290 458334 528390 458434
rect 528514 458334 528592 458434
rect 528592 458334 528614 458434
rect 527618 458110 527718 458210
rect 527842 458110 527942 458210
rect 528066 458110 528166 458210
rect 528290 458110 528390 458210
rect 528514 458110 528592 458210
rect 528592 458110 528614 458210
rect 527618 457886 527718 457986
rect 527842 457886 527942 457986
rect 528066 457886 528166 457986
rect 528290 457886 528390 457986
rect 528514 457886 528592 457986
rect 528592 457886 528614 457986
rect 527618 457662 527718 457762
rect 527842 457662 527942 457762
rect 528066 457662 528166 457762
rect 528290 457662 528390 457762
rect 528514 457662 528592 457762
rect 528592 457662 528614 457762
rect 527618 457438 527718 457538
rect 527842 457438 527942 457538
rect 528066 457438 528166 457538
rect 528290 457438 528390 457538
rect 528514 457438 528592 457538
rect 528592 457438 528614 457538
rect 527618 457214 527718 457314
rect 527842 457214 527942 457314
rect 528066 457214 528166 457314
rect 528290 457214 528390 457314
rect 528514 457214 528592 457314
rect 528592 457214 528614 457314
rect 562190 455178 562252 455212
rect 562252 455178 567482 455212
rect 567482 455178 567544 455212
rect 562156 454073 562190 455055
rect 562270 454112 562304 455088
rect 562528 454112 562562 455088
rect 562786 454112 562820 455088
rect 563044 454112 563078 455088
rect 563302 454112 563336 455088
rect 563560 454112 563594 455088
rect 563818 454112 563852 455088
rect 564076 454112 564110 455088
rect 564334 454112 564368 455088
rect 564592 454112 564626 455088
rect 564850 454112 564884 455088
rect 565108 454112 565142 455088
rect 565366 454112 565400 455088
rect 565624 454112 565658 455088
rect 565882 454112 565916 455088
rect 566140 454112 566174 455088
rect 566398 454112 566432 455088
rect 566656 454112 566690 455088
rect 566914 454112 566948 455088
rect 567172 454112 567206 455088
rect 567430 454112 567464 455088
rect 567544 454073 567578 455055
rect 562374 454019 562458 454053
rect 562632 454019 562716 454053
rect 562890 454019 562974 454053
rect 563148 454019 563232 454053
rect 563406 454019 563490 454053
rect 563664 454019 563748 454053
rect 563922 454019 564006 454053
rect 564180 454019 564264 454053
rect 564438 454019 564522 454053
rect 564696 454019 564780 454053
rect 564954 454019 565038 454053
rect 565212 454019 565296 454053
rect 565470 454019 565554 454053
rect 565728 454019 565812 454053
rect 565986 454019 566070 454053
rect 566244 454019 566328 454053
rect 566502 454019 566586 454053
rect 566760 454019 566844 454053
rect 567018 454019 567102 454053
rect 567276 454019 567360 454053
rect 572350 455212 572412 455246
rect 572412 455212 577642 455246
rect 577642 455212 577704 455246
rect 572316 454116 572350 455090
rect 572430 454146 572464 455122
rect 572688 454146 572722 455122
rect 572946 454146 572980 455122
rect 573204 454146 573238 455122
rect 573462 454146 573496 455122
rect 573720 454146 573754 455122
rect 573978 454146 574012 455122
rect 574236 454146 574270 455122
rect 574494 454146 574528 455122
rect 574752 454146 574786 455122
rect 575010 454146 575044 455122
rect 575268 454146 575302 455122
rect 575526 454146 575560 455122
rect 575784 454146 575818 455122
rect 576042 454146 576076 455122
rect 576300 454146 576334 455122
rect 576558 454146 576592 455122
rect 576816 454146 576850 455122
rect 577074 454146 577108 455122
rect 577332 454146 577366 455122
rect 577590 454146 577624 455122
rect 577704 454116 577738 455090
rect 572534 454062 572618 454096
rect 572792 454062 572876 454096
rect 573050 454062 573134 454096
rect 573308 454062 573392 454096
rect 573566 454062 573650 454096
rect 573824 454062 573908 454096
rect 574082 454062 574166 454096
rect 574340 454062 574424 454096
rect 574598 454062 574682 454096
rect 574856 454062 574940 454096
rect 575114 454062 575198 454096
rect 575372 454062 575456 454096
rect 575630 454062 575714 454096
rect 575888 454062 575972 454096
rect 576146 454062 576230 454096
rect 576404 454062 576488 454096
rect 576662 454062 576746 454096
rect 576920 454062 577004 454096
rect 577178 454062 577262 454096
rect 577436 454062 577520 454096
rect 527638 437440 527738 437540
rect 527862 437440 527962 437540
rect 528086 437440 528186 437540
rect 528310 437440 528410 437540
rect 528534 437440 528592 437540
rect 528592 437440 528634 437540
rect 527638 437216 527738 437316
rect 527862 437216 527962 437316
rect 528086 437216 528186 437316
rect 528310 437216 528410 437316
rect 528534 437216 528592 437316
rect 528592 437216 528634 437316
rect 527638 436992 527738 437092
rect 527862 436992 527962 437092
rect 528086 436992 528186 437092
rect 528310 436992 528410 437092
rect 528534 436992 528592 437092
rect 528592 436992 528634 437092
rect 527638 436768 527738 436868
rect 527862 436768 527962 436868
rect 528086 436768 528186 436868
rect 528310 436768 528410 436868
rect 528534 436768 528592 436868
rect 528592 436768 528634 436868
rect 527638 436544 527738 436644
rect 527862 436544 527962 436644
rect 528086 436544 528186 436644
rect 528310 436544 528410 436644
rect 528534 436544 528592 436644
rect 528592 436544 528634 436644
rect 527638 436320 527738 436420
rect 527862 436320 527962 436420
rect 528086 436320 528186 436420
rect 528310 436320 528410 436420
rect 528534 436320 528592 436420
rect 528592 436320 528634 436420
rect 527638 436096 527738 436196
rect 527862 436096 527962 436196
rect 528086 436096 528186 436196
rect 528310 436096 528410 436196
rect 528534 436096 528592 436196
rect 528592 436096 528634 436196
rect 527638 435872 527738 435972
rect 527862 435872 527962 435972
rect 528086 435872 528186 435972
rect 528310 435872 528410 435972
rect 528534 435872 528592 435972
rect 528592 435872 528634 435972
rect 527638 435648 527738 435748
rect 527862 435648 527962 435748
rect 528086 435648 528186 435748
rect 528310 435648 528410 435748
rect 528534 435648 528592 435748
rect 528592 435648 528634 435748
rect 527638 435424 527738 435524
rect 527862 435424 527962 435524
rect 528086 435424 528186 435524
rect 528310 435424 528410 435524
rect 528534 435424 528592 435524
rect 528592 435424 528634 435524
rect 527638 435200 527738 435300
rect 527862 435200 527962 435300
rect 528086 435200 528186 435300
rect 528310 435200 528410 435300
rect 528534 435200 528592 435300
rect 528592 435200 528634 435300
rect 527638 434976 527738 435076
rect 527862 434976 527962 435076
rect 528086 434976 528186 435076
rect 528310 434976 528410 435076
rect 528534 434976 528592 435076
rect 528592 434976 528634 435076
rect 527638 434752 527738 434852
rect 527862 434752 527962 434852
rect 528086 434752 528186 434852
rect 528310 434752 528410 434852
rect 528534 434752 528592 434852
rect 528592 434752 528634 434852
rect 527638 434528 527738 434628
rect 527862 434528 527962 434628
rect 528086 434528 528186 434628
rect 528310 434528 528410 434628
rect 528534 434528 528592 434628
rect 528592 434528 528634 434628
rect 527638 434304 527738 434404
rect 527862 434304 527962 434404
rect 528086 434304 528186 434404
rect 528310 434304 528410 434404
rect 528534 434304 528592 434404
rect 528592 434304 528634 434404
rect 527638 434080 527738 434180
rect 527862 434080 527962 434180
rect 528086 434080 528186 434180
rect 528310 434080 528410 434180
rect 528534 434080 528592 434180
rect 528592 434080 528634 434180
rect 527638 433856 527738 433956
rect 527862 433856 527962 433956
rect 528086 433856 528186 433956
rect 528310 433856 528410 433956
rect 528534 433856 528592 433956
rect 528592 433856 528634 433956
rect 527638 433632 527738 433732
rect 527862 433632 527962 433732
rect 528086 433632 528186 433732
rect 528310 433632 528410 433732
rect 528534 433632 528592 433732
rect 528592 433632 528634 433732
rect 527638 433408 527738 433508
rect 527862 433408 527962 433508
rect 528086 433408 528186 433508
rect 528310 433408 528410 433508
rect 528534 433408 528592 433508
rect 528592 433408 528634 433508
rect 527638 433184 527738 433284
rect 527862 433184 527962 433284
rect 528086 433184 528186 433284
rect 528310 433184 528410 433284
rect 528534 433184 528592 433284
rect 528592 433184 528634 433284
rect 527638 432960 527738 433060
rect 527862 432960 527962 433060
rect 528086 432960 528186 433060
rect 528310 432960 528410 433060
rect 528534 432960 528592 433060
rect 528592 432960 528634 433060
rect 527638 432736 527738 432836
rect 527862 432736 527962 432836
rect 528086 432736 528186 432836
rect 528310 432736 528410 432836
rect 528534 432736 528592 432836
rect 528592 432736 528634 432836
rect 527638 432512 527738 432612
rect 527862 432512 527962 432612
rect 528086 432512 528186 432612
rect 528310 432512 528410 432612
rect 528534 432512 528592 432612
rect 528592 432512 528634 432612
rect 527638 432288 527738 432388
rect 527862 432288 527962 432388
rect 528086 432288 528186 432388
rect 528310 432288 528410 432388
rect 528534 432288 528592 432388
rect 528592 432288 528634 432388
rect 527638 432064 527738 432164
rect 527862 432064 527962 432164
rect 528086 432064 528186 432164
rect 528310 432064 528410 432164
rect 528534 432064 528592 432164
rect 528592 432064 528634 432164
rect 527638 431840 527738 431940
rect 527862 431840 527962 431940
rect 528086 431840 528186 431940
rect 528310 431840 528410 431940
rect 528534 431840 528592 431940
rect 528592 431840 528634 431940
rect 527638 431616 527738 431716
rect 527862 431616 527962 431716
rect 528086 431616 528186 431716
rect 528310 431616 528410 431716
rect 528534 431616 528592 431716
rect 528592 431616 528634 431716
rect 527638 431392 527738 431492
rect 527862 431392 527962 431492
rect 528086 431392 528186 431492
rect 528310 431392 528410 431492
rect 528534 431392 528592 431492
rect 528592 431392 528634 431492
rect 527638 431168 527738 431268
rect 527862 431168 527962 431268
rect 528086 431168 528186 431268
rect 528310 431168 528410 431268
rect 528534 431168 528592 431268
rect 528592 431168 528634 431268
rect 503920 430702 504020 430802
rect 504144 430702 504244 430802
rect 504368 430702 504468 430802
rect 504592 430702 504692 430802
rect 504816 430702 504916 430802
rect 505040 430702 505140 430802
rect 505264 430702 505364 430802
rect 505488 430702 505588 430802
rect 505712 430702 505812 430802
rect 505936 430702 506036 430802
rect 506160 430702 506260 430802
rect 506384 430702 506484 430802
rect 506608 430702 506708 430802
rect 506832 430702 506932 430802
rect 507056 430702 507156 430802
rect 507280 430702 507380 430802
rect 507504 430702 507604 430802
rect 507728 430702 507828 430802
rect 507952 430702 508052 430802
rect 508176 430702 508276 430802
rect 508400 430702 508500 430802
rect 508624 430702 508724 430802
rect 508848 430702 508948 430802
rect 509072 430702 509172 430802
rect 509296 430702 509396 430802
rect 509520 430702 509620 430802
rect 509744 430702 509844 430802
rect 509968 430702 510068 430802
rect 510192 430702 510292 430802
rect 510416 430702 510516 430802
rect 517320 430702 517420 430802
rect 517544 430702 517644 430802
rect 517768 430702 517868 430802
rect 517992 430702 518092 430802
rect 518216 430702 518316 430802
rect 518440 430702 518540 430802
rect 518664 430702 518764 430802
rect 518888 430702 518988 430802
rect 519112 430702 519212 430802
rect 519336 430702 519436 430802
rect 519560 430702 519660 430802
rect 519784 430702 519884 430802
rect 520008 430702 520108 430802
rect 520232 430702 520332 430802
rect 520456 430702 520556 430802
rect 520680 430702 520780 430802
rect 520904 430702 521004 430802
rect 521128 430702 521228 430802
rect 521352 430702 521452 430802
rect 521576 430702 521676 430802
rect 521800 430702 521900 430802
rect 522024 430702 522124 430802
rect 522248 430702 522348 430802
rect 522472 430702 522572 430802
rect 522696 430702 522796 430802
rect 522920 430702 523020 430802
rect 523144 430702 523244 430802
rect 523368 430702 523468 430802
rect 523592 430702 523692 430802
rect 523816 430702 523916 430802
rect 503920 430478 504020 430578
rect 504144 430478 504244 430578
rect 504368 430478 504468 430578
rect 504592 430478 504692 430578
rect 504816 430478 504916 430578
rect 505040 430478 505140 430578
rect 505264 430478 505364 430578
rect 505488 430478 505588 430578
rect 505712 430478 505812 430578
rect 505936 430478 506036 430578
rect 506160 430478 506260 430578
rect 506384 430478 506484 430578
rect 506608 430478 506708 430578
rect 506832 430478 506932 430578
rect 507056 430478 507156 430578
rect 507280 430478 507380 430578
rect 507504 430478 507604 430578
rect 507728 430478 507828 430578
rect 507952 430478 508052 430578
rect 508176 430478 508276 430578
rect 508400 430478 508500 430578
rect 508624 430478 508724 430578
rect 508848 430478 508948 430578
rect 509072 430478 509172 430578
rect 509296 430478 509396 430578
rect 509520 430478 509620 430578
rect 509744 430478 509844 430578
rect 509968 430478 510068 430578
rect 510192 430478 510292 430578
rect 510416 430478 510516 430578
rect 517320 430478 517420 430578
rect 517544 430478 517644 430578
rect 517768 430478 517868 430578
rect 517992 430478 518092 430578
rect 518216 430478 518316 430578
rect 518440 430478 518540 430578
rect 518664 430478 518764 430578
rect 518888 430478 518988 430578
rect 519112 430478 519212 430578
rect 519336 430478 519436 430578
rect 519560 430478 519660 430578
rect 519784 430478 519884 430578
rect 520008 430478 520108 430578
rect 520232 430478 520332 430578
rect 520456 430478 520556 430578
rect 520680 430478 520780 430578
rect 520904 430478 521004 430578
rect 521128 430478 521228 430578
rect 521352 430478 521452 430578
rect 521576 430478 521676 430578
rect 521800 430478 521900 430578
rect 522024 430478 522124 430578
rect 522248 430478 522348 430578
rect 522472 430478 522572 430578
rect 522696 430478 522796 430578
rect 522920 430478 523020 430578
rect 523144 430478 523244 430578
rect 523368 430478 523468 430578
rect 523592 430478 523692 430578
rect 523816 430478 523916 430578
rect 503920 430254 504020 430354
rect 504144 430254 504244 430354
rect 504368 430254 504468 430354
rect 504592 430254 504692 430354
rect 504816 430254 504916 430354
rect 505040 430254 505140 430354
rect 505264 430254 505364 430354
rect 505488 430254 505588 430354
rect 505712 430254 505812 430354
rect 505936 430254 506036 430354
rect 506160 430254 506260 430354
rect 506384 430254 506484 430354
rect 506608 430254 506708 430354
rect 506832 430254 506932 430354
rect 507056 430254 507156 430354
rect 507280 430254 507380 430354
rect 507504 430254 507604 430354
rect 507728 430254 507828 430354
rect 507952 430254 508052 430354
rect 508176 430254 508276 430354
rect 508400 430254 508500 430354
rect 508624 430254 508724 430354
rect 508848 430254 508948 430354
rect 509072 430254 509172 430354
rect 509296 430254 509396 430354
rect 509520 430254 509620 430354
rect 509744 430254 509844 430354
rect 509968 430254 510068 430354
rect 510192 430254 510292 430354
rect 510416 430254 510516 430354
rect 517320 430254 517420 430354
rect 517544 430254 517644 430354
rect 517768 430254 517868 430354
rect 517992 430254 518092 430354
rect 518216 430254 518316 430354
rect 518440 430254 518540 430354
rect 518664 430254 518764 430354
rect 518888 430254 518988 430354
rect 519112 430254 519212 430354
rect 519336 430254 519436 430354
rect 519560 430254 519660 430354
rect 519784 430254 519884 430354
rect 520008 430254 520108 430354
rect 520232 430254 520332 430354
rect 520456 430254 520556 430354
rect 520680 430254 520780 430354
rect 520904 430254 521004 430354
rect 521128 430254 521228 430354
rect 521352 430254 521452 430354
rect 521576 430254 521676 430354
rect 521800 430254 521900 430354
rect 522024 430254 522124 430354
rect 522248 430254 522348 430354
rect 522472 430254 522572 430354
rect 522696 430254 522796 430354
rect 522920 430254 523020 430354
rect 523144 430254 523244 430354
rect 523368 430254 523468 430354
rect 523592 430254 523692 430354
rect 523816 430254 523916 430354
rect 503920 430044 504020 430130
rect 504144 430044 504244 430130
rect 504368 430044 504468 430130
rect 504592 430044 504692 430130
rect 504816 430044 504916 430130
rect 505040 430044 505140 430130
rect 505264 430044 505364 430130
rect 505488 430044 505588 430130
rect 505712 430044 505812 430130
rect 505936 430044 506036 430130
rect 506160 430044 506260 430130
rect 506384 430044 506484 430130
rect 506608 430044 506708 430130
rect 506832 430044 506932 430130
rect 507056 430044 507156 430130
rect 507280 430044 507380 430130
rect 507504 430044 507604 430130
rect 507728 430044 507828 430130
rect 507952 430044 508052 430130
rect 508176 430044 508276 430130
rect 508400 430044 508500 430130
rect 508624 430044 508724 430130
rect 508848 430044 508948 430130
rect 509072 430044 509172 430130
rect 509296 430044 509396 430130
rect 509520 430044 509620 430130
rect 509744 430044 509844 430130
rect 509968 430044 510068 430130
rect 510192 430044 510292 430130
rect 510416 430044 510516 430130
rect 517320 430044 517420 430130
rect 517544 430044 517644 430130
rect 517768 430044 517868 430130
rect 517992 430044 518092 430130
rect 518216 430044 518316 430130
rect 518440 430044 518540 430130
rect 518664 430044 518764 430130
rect 518888 430044 518988 430130
rect 519112 430044 519212 430130
rect 519336 430044 519436 430130
rect 519560 430044 519660 430130
rect 519784 430044 519884 430130
rect 520008 430044 520108 430130
rect 520232 430044 520332 430130
rect 520456 430044 520556 430130
rect 520680 430044 520780 430130
rect 520904 430044 521004 430130
rect 521128 430044 521228 430130
rect 521352 430044 521452 430130
rect 521576 430044 521676 430130
rect 521800 430044 521900 430130
rect 522024 430044 522124 430130
rect 522248 430044 522348 430130
rect 522472 430044 522572 430130
rect 522696 430044 522796 430130
rect 522920 430044 523020 430130
rect 523144 430044 523244 430130
rect 523368 430044 523468 430130
rect 523592 430044 523692 430130
rect 523816 430044 523916 430130
rect 527638 430944 527738 431044
rect 527862 430944 527962 431044
rect 528086 430944 528186 431044
rect 528310 430944 528410 431044
rect 528534 430944 528592 431044
rect 528592 430944 528634 431044
rect 503920 430030 504020 430044
rect 504144 430030 504244 430044
rect 504368 430030 504468 430044
rect 504592 430030 504692 430044
rect 504816 430030 504916 430044
rect 505040 430030 505140 430044
rect 505264 430030 505364 430044
rect 505488 430030 505588 430044
rect 505712 430030 505812 430044
rect 505936 430030 506036 430044
rect 506160 430030 506260 430044
rect 506384 430030 506484 430044
rect 506608 430030 506708 430044
rect 506832 430030 506932 430044
rect 507056 430030 507156 430044
rect 507280 430030 507380 430044
rect 507504 430030 507604 430044
rect 507728 430030 507828 430044
rect 507952 430030 508052 430044
rect 508176 430030 508276 430044
rect 508400 430030 508500 430044
rect 508624 430030 508724 430044
rect 508848 430030 508948 430044
rect 509072 430030 509172 430044
rect 509296 430030 509396 430044
rect 509520 430030 509620 430044
rect 509744 430030 509844 430044
rect 509968 430030 510068 430044
rect 510192 430030 510292 430044
rect 510416 430030 510516 430044
rect 517320 430030 517420 430044
rect 517544 430030 517644 430044
rect 517768 430030 517868 430044
rect 517992 430030 518092 430044
rect 518216 430030 518316 430044
rect 518440 430030 518540 430044
rect 518664 430030 518764 430044
rect 518888 430030 518988 430044
rect 519112 430030 519212 430044
rect 519336 430030 519436 430044
rect 519560 430030 519660 430044
rect 519784 430030 519884 430044
rect 520008 430030 520108 430044
rect 520232 430030 520332 430044
rect 520456 430030 520556 430044
rect 520680 430030 520780 430044
rect 520904 430030 521004 430044
rect 521128 430030 521228 430044
rect 521352 430030 521452 430044
rect 521576 430030 521676 430044
rect 521800 430030 521900 430044
rect 522024 430030 522124 430044
rect 522248 430030 522348 430044
rect 522472 430030 522572 430044
rect 522696 430030 522796 430044
rect 522920 430030 523020 430044
rect 523144 430030 523244 430044
rect 523368 430030 523468 430044
rect 523592 430030 523692 430044
rect 523816 430030 523916 430044
<< metal1 >>
rect 562150 495742 567584 495775
rect 562150 495662 562480 495742
rect 562560 495662 562640 495742
rect 562720 495662 562800 495742
rect 562880 495662 562960 495742
rect 563040 495662 563120 495742
rect 563200 495662 563280 495742
rect 563360 495662 563440 495742
rect 563520 495662 563600 495742
rect 563680 495662 563760 495742
rect 563840 495662 563920 495742
rect 564000 495662 564080 495742
rect 564160 495662 564240 495742
rect 564320 495662 564400 495742
rect 564480 495662 564560 495742
rect 564640 495662 564720 495742
rect 564800 495662 564880 495742
rect 564960 495662 565040 495742
rect 565120 495662 565200 495742
rect 565280 495662 565360 495742
rect 565440 495662 565520 495742
rect 565600 495662 565680 495742
rect 565760 495662 565840 495742
rect 565920 495662 566000 495742
rect 566080 495662 566160 495742
rect 566240 495662 566320 495742
rect 566400 495662 566480 495742
rect 566560 495662 566640 495742
rect 566720 495662 566800 495742
rect 566880 495662 566960 495742
rect 567040 495662 567120 495742
rect 567200 495662 567280 495742
rect 567360 495662 567584 495742
rect 562150 495582 567584 495662
rect 562150 495514 562480 495582
rect 562560 495514 562640 495582
rect 562720 495514 562800 495582
rect 562880 495514 562960 495582
rect 563040 495514 563120 495582
rect 563200 495514 563280 495582
rect 563360 495514 563440 495582
rect 563520 495514 563600 495582
rect 563680 495514 563760 495582
rect 563840 495514 563920 495582
rect 564000 495514 564080 495582
rect 564160 495514 564240 495582
rect 564320 495514 564400 495582
rect 564480 495514 564560 495582
rect 564640 495514 564720 495582
rect 564800 495514 564880 495582
rect 564960 495514 565040 495582
rect 565120 495514 565200 495582
rect 565280 495514 565360 495582
rect 565440 495514 565520 495582
rect 565600 495514 565680 495582
rect 565760 495514 565840 495582
rect 565920 495514 566000 495582
rect 566080 495514 566160 495582
rect 566240 495514 566320 495582
rect 566400 495514 566480 495582
rect 566560 495514 566640 495582
rect 566720 495514 566800 495582
rect 566880 495514 566960 495582
rect 567040 495514 567120 495582
rect 567200 495514 567280 495582
rect 567360 495514 567584 495582
rect 562150 495480 562190 495514
rect 567544 495480 567584 495514
rect 562150 495474 567584 495480
rect 562150 495357 562196 495474
rect 562150 494375 562156 495357
rect 562190 494375 562196 495357
rect 562150 494363 562196 494375
rect 562264 495390 562310 495402
rect 562264 494414 562270 495390
rect 562304 494414 562310 495390
rect 562264 494277 562310 494414
rect 562522 495390 562568 495474
rect 562522 494414 562528 495390
rect 562562 494414 562568 495390
rect 562522 494402 562568 494414
rect 562780 495390 562826 495402
rect 562780 494414 562786 495390
rect 562820 494414 562826 495390
rect 562362 494355 562470 494361
rect 562362 494321 562374 494355
rect 562458 494321 562470 494355
rect 562362 494315 562470 494321
rect 562620 494355 562728 494361
rect 562620 494321 562632 494355
rect 562716 494321 562728 494355
rect 562620 494315 562728 494321
rect 562780 494277 562826 494414
rect 563038 495390 563084 495474
rect 563038 494414 563044 495390
rect 563078 494414 563084 495390
rect 563038 494402 563084 494414
rect 563296 495390 563342 495402
rect 563296 494414 563302 495390
rect 563336 494414 563342 495390
rect 562878 494355 562986 494361
rect 562878 494321 562890 494355
rect 562974 494321 562986 494355
rect 562878 494315 562986 494321
rect 563136 494355 563244 494361
rect 563136 494321 563148 494355
rect 563232 494321 563244 494355
rect 563136 494315 563244 494321
rect 563296 494277 563342 494414
rect 563554 495390 563600 495474
rect 563554 494414 563560 495390
rect 563594 494414 563600 495390
rect 563554 494402 563600 494414
rect 563812 495390 563858 495402
rect 563812 494414 563818 495390
rect 563852 494414 563858 495390
rect 563394 494355 563502 494361
rect 563394 494321 563406 494355
rect 563490 494321 563502 494355
rect 563394 494315 563502 494321
rect 563652 494355 563760 494361
rect 563652 494321 563664 494355
rect 563748 494321 563760 494355
rect 563652 494315 563760 494321
rect 563812 494277 563858 494414
rect 564070 495390 564116 495474
rect 564070 494414 564076 495390
rect 564110 494414 564116 495390
rect 564070 494402 564116 494414
rect 564328 495390 564374 495402
rect 564328 494414 564334 495390
rect 564368 494414 564374 495390
rect 563910 494355 564018 494361
rect 563910 494321 563922 494355
rect 564006 494321 564018 494355
rect 563910 494315 564018 494321
rect 564168 494355 564276 494361
rect 564168 494321 564180 494355
rect 564264 494321 564276 494355
rect 564168 494315 564276 494321
rect 564328 494277 564374 494414
rect 564586 495390 564632 495474
rect 564586 494414 564592 495390
rect 564626 494414 564632 495390
rect 564586 494402 564632 494414
rect 564844 495390 564890 495402
rect 564844 494414 564850 495390
rect 564884 494414 564890 495390
rect 564426 494355 564534 494361
rect 564426 494321 564438 494355
rect 564522 494321 564534 494355
rect 564426 494315 564534 494321
rect 564684 494355 564792 494361
rect 564684 494321 564696 494355
rect 564780 494321 564792 494355
rect 564684 494315 564792 494321
rect 564844 494277 564890 494414
rect 565102 495390 565148 495474
rect 565102 494414 565108 495390
rect 565142 494414 565148 495390
rect 565102 494402 565148 494414
rect 565360 495390 565406 495402
rect 565360 494414 565366 495390
rect 565400 494414 565406 495390
rect 564942 494355 565050 494361
rect 564942 494321 564954 494355
rect 565038 494321 565050 494355
rect 564942 494315 565050 494321
rect 565200 494355 565308 494361
rect 565200 494321 565212 494355
rect 565296 494321 565308 494355
rect 565200 494315 565308 494321
rect 565360 494277 565406 494414
rect 565618 495390 565664 495474
rect 565618 494414 565624 495390
rect 565658 494414 565664 495390
rect 565618 494402 565664 494414
rect 565876 495390 565922 495402
rect 565876 494414 565882 495390
rect 565916 494414 565922 495390
rect 565458 494355 565566 494361
rect 565458 494321 565470 494355
rect 565554 494321 565566 494355
rect 565458 494315 565566 494321
rect 565716 494355 565824 494361
rect 565716 494321 565728 494355
rect 565812 494321 565824 494355
rect 565716 494315 565824 494321
rect 565876 494277 565922 494414
rect 566134 495390 566180 495474
rect 566134 494414 566140 495390
rect 566174 494414 566180 495390
rect 566134 494402 566180 494414
rect 566392 495390 566438 495402
rect 566392 494414 566398 495390
rect 566432 494414 566438 495390
rect 565974 494355 566082 494361
rect 565974 494321 565986 494355
rect 566070 494321 566082 494355
rect 565974 494315 566082 494321
rect 566232 494355 566340 494361
rect 566232 494321 566244 494355
rect 566328 494321 566340 494355
rect 566232 494315 566340 494321
rect 566392 494277 566438 494414
rect 566650 495390 566696 495474
rect 566650 494414 566656 495390
rect 566690 494414 566696 495390
rect 566650 494402 566696 494414
rect 566908 495390 566954 495402
rect 566908 494414 566914 495390
rect 566948 494414 566954 495390
rect 566490 494355 566598 494361
rect 566490 494321 566502 494355
rect 566586 494321 566598 494355
rect 566490 494315 566598 494321
rect 566748 494355 566856 494361
rect 566748 494321 566760 494355
rect 566844 494321 566856 494355
rect 566748 494315 566856 494321
rect 566908 494277 566954 494414
rect 567166 495390 567212 495474
rect 567166 494414 567172 495390
rect 567206 494414 567212 495390
rect 567166 494402 567212 494414
rect 567424 495390 567470 495402
rect 567424 494414 567430 495390
rect 567464 494414 567470 495390
rect 567006 494355 567114 494361
rect 567006 494321 567018 494355
rect 567102 494321 567114 494355
rect 567006 494315 567114 494321
rect 567264 494355 567372 494361
rect 567264 494321 567276 494355
rect 567360 494321 567372 494355
rect 567264 494315 567372 494321
rect 567424 494277 567470 494414
rect 567538 495357 567584 495474
rect 567538 494375 567544 495357
rect 567578 494375 567584 495357
rect 572310 495742 577744 495775
rect 572310 495662 572640 495742
rect 572720 495662 572800 495742
rect 572880 495662 572960 495742
rect 573040 495662 573120 495742
rect 573200 495662 573280 495742
rect 573360 495662 573440 495742
rect 573520 495662 573600 495742
rect 573680 495662 573760 495742
rect 573840 495662 573920 495742
rect 574000 495662 574080 495742
rect 574160 495662 574240 495742
rect 574320 495662 574400 495742
rect 574480 495662 574560 495742
rect 574640 495662 574720 495742
rect 574800 495662 574880 495742
rect 574960 495662 575040 495742
rect 575120 495662 575200 495742
rect 575280 495662 575360 495742
rect 575440 495662 575520 495742
rect 575600 495662 575680 495742
rect 575760 495662 575840 495742
rect 575920 495662 576000 495742
rect 576080 495662 576160 495742
rect 576240 495662 576320 495742
rect 576400 495662 576480 495742
rect 576560 495662 576640 495742
rect 576720 495662 576800 495742
rect 576880 495662 576960 495742
rect 577040 495662 577120 495742
rect 577200 495662 577280 495742
rect 577360 495662 577440 495742
rect 577520 495662 577744 495742
rect 572310 495582 577744 495662
rect 572310 495548 572640 495582
rect 572720 495548 572800 495582
rect 572880 495548 572960 495582
rect 573040 495548 573120 495582
rect 573200 495548 573280 495582
rect 573360 495548 573440 495582
rect 573520 495548 573600 495582
rect 573680 495548 573760 495582
rect 573840 495548 573920 495582
rect 574000 495548 574080 495582
rect 574160 495548 574240 495582
rect 574320 495548 574400 495582
rect 574480 495548 574560 495582
rect 574640 495548 574720 495582
rect 574800 495548 574880 495582
rect 574960 495548 575040 495582
rect 575120 495548 575200 495582
rect 575280 495548 575360 495582
rect 575440 495548 575520 495582
rect 575600 495548 575680 495582
rect 575760 495548 575840 495582
rect 575920 495548 576000 495582
rect 576080 495548 576160 495582
rect 576240 495548 576320 495582
rect 576400 495548 576480 495582
rect 576560 495548 576640 495582
rect 576720 495548 576800 495582
rect 576880 495548 576960 495582
rect 577040 495548 577120 495582
rect 577200 495548 577280 495582
rect 577360 495548 577440 495582
rect 577520 495548 577744 495582
rect 572310 495514 572350 495548
rect 577704 495514 577744 495548
rect 572310 495502 572640 495514
rect 572720 495502 572800 495514
rect 572880 495502 572960 495514
rect 573040 495502 573120 495514
rect 573200 495502 573280 495514
rect 573360 495502 573440 495514
rect 573520 495502 573600 495514
rect 573680 495502 573760 495514
rect 573840 495502 573920 495514
rect 574000 495502 574080 495514
rect 574160 495502 574240 495514
rect 574320 495502 574400 495514
rect 574480 495502 574560 495514
rect 574640 495502 574720 495514
rect 574800 495502 574880 495514
rect 574960 495502 575040 495514
rect 575120 495502 575200 495514
rect 575280 495502 575360 495514
rect 575440 495502 575520 495514
rect 575600 495502 575680 495514
rect 575760 495502 575840 495514
rect 575920 495502 576000 495514
rect 576080 495502 576160 495514
rect 576240 495502 576320 495514
rect 576400 495502 576480 495514
rect 576560 495502 576640 495514
rect 576720 495502 576800 495514
rect 576880 495502 576960 495514
rect 577040 495502 577120 495514
rect 577200 495502 577280 495514
rect 577360 495502 577440 495514
rect 577520 495502 577744 495514
rect 572310 495474 577744 495502
rect 572310 495392 572356 495474
rect 572688 495436 572722 495474
rect 573204 495436 573238 495474
rect 573720 495436 573754 495474
rect 574236 495436 574270 495474
rect 574752 495436 574786 495474
rect 575268 495436 575302 495474
rect 575784 495436 575818 495474
rect 576300 495436 576334 495474
rect 576816 495436 576850 495474
rect 577332 495436 577366 495474
rect 572310 494418 572316 495392
rect 572350 494418 572356 495392
rect 572310 494406 572356 494418
rect 572424 495424 572470 495436
rect 572424 494448 572430 495424
rect 572464 494448 572470 495424
rect 567538 494363 567584 494375
rect 572424 494292 572470 494448
rect 572682 495424 572728 495436
rect 572682 494448 572688 495424
rect 572722 494448 572728 495424
rect 572682 494436 572728 494448
rect 572940 495424 572986 495436
rect 572940 494448 572946 495424
rect 572980 494448 572986 495424
rect 572522 494398 572630 494404
rect 572522 494364 572534 494398
rect 572618 494364 572630 494398
rect 572522 494358 572630 494364
rect 572780 494398 572888 494404
rect 572780 494364 572792 494398
rect 572876 494364 572888 494398
rect 572780 494358 572888 494364
rect 572940 494292 572986 494448
rect 573198 495424 573244 495436
rect 573198 494448 573204 495424
rect 573238 494448 573244 495424
rect 573198 494436 573244 494448
rect 573456 495424 573502 495436
rect 573456 494448 573462 495424
rect 573496 494448 573502 495424
rect 573038 494398 573146 494404
rect 573038 494364 573050 494398
rect 573134 494364 573146 494398
rect 573038 494358 573146 494364
rect 573296 494398 573404 494404
rect 573296 494364 573308 494398
rect 573392 494364 573404 494398
rect 573296 494358 573404 494364
rect 573456 494292 573502 494448
rect 573714 495424 573760 495436
rect 573714 494448 573720 495424
rect 573754 494448 573760 495424
rect 573714 494436 573760 494448
rect 573972 495424 574018 495436
rect 573972 494448 573978 495424
rect 574012 494448 574018 495424
rect 573554 494398 573662 494404
rect 573554 494364 573566 494398
rect 573650 494364 573662 494398
rect 573554 494358 573662 494364
rect 573812 494398 573920 494404
rect 573812 494364 573824 494398
rect 573908 494364 573920 494398
rect 573812 494358 573920 494364
rect 573972 494292 574018 494448
rect 574230 495424 574276 495436
rect 574230 494448 574236 495424
rect 574270 494448 574276 495424
rect 574230 494436 574276 494448
rect 574488 495424 574534 495436
rect 574488 494448 574494 495424
rect 574528 494448 574534 495424
rect 574070 494398 574178 494404
rect 574070 494364 574082 494398
rect 574166 494364 574178 494398
rect 574070 494358 574178 494364
rect 574328 494398 574436 494404
rect 574328 494364 574340 494398
rect 574424 494364 574436 494398
rect 574328 494358 574436 494364
rect 574488 494292 574534 494448
rect 574746 495424 574792 495436
rect 574746 494448 574752 495424
rect 574786 494448 574792 495424
rect 574746 494436 574792 494448
rect 575004 495424 575050 495436
rect 575004 494448 575010 495424
rect 575044 494448 575050 495424
rect 574586 494398 574694 494404
rect 574586 494364 574598 494398
rect 574682 494364 574694 494398
rect 574586 494358 574694 494364
rect 574844 494398 574952 494404
rect 574844 494364 574856 494398
rect 574940 494364 574952 494398
rect 574844 494358 574952 494364
rect 575004 494292 575050 494448
rect 575262 495424 575308 495436
rect 575262 494448 575268 495424
rect 575302 494448 575308 495424
rect 575262 494436 575308 494448
rect 575520 495424 575566 495436
rect 575520 494448 575526 495424
rect 575560 494448 575566 495424
rect 575102 494398 575210 494404
rect 575102 494364 575114 494398
rect 575198 494364 575210 494398
rect 575102 494358 575210 494364
rect 575360 494398 575468 494404
rect 575360 494364 575372 494398
rect 575456 494364 575468 494398
rect 575360 494358 575468 494364
rect 575520 494292 575566 494448
rect 575778 495424 575824 495436
rect 575778 494448 575784 495424
rect 575818 494448 575824 495424
rect 575778 494436 575824 494448
rect 576036 495424 576082 495436
rect 576036 494448 576042 495424
rect 576076 494448 576082 495424
rect 575618 494398 575726 494404
rect 575618 494364 575630 494398
rect 575714 494364 575726 494398
rect 575618 494358 575726 494364
rect 575876 494398 575984 494404
rect 575876 494364 575888 494398
rect 575972 494364 575984 494398
rect 575876 494358 575984 494364
rect 576036 494292 576082 494448
rect 576294 495424 576340 495436
rect 576294 494448 576300 495424
rect 576334 494448 576340 495424
rect 576294 494436 576340 494448
rect 576552 495424 576598 495436
rect 576552 494448 576558 495424
rect 576592 494448 576598 495424
rect 576134 494398 576242 494404
rect 576134 494364 576146 494398
rect 576230 494364 576242 494398
rect 576134 494358 576242 494364
rect 576392 494398 576500 494404
rect 576392 494364 576404 494398
rect 576488 494364 576500 494398
rect 576392 494358 576500 494364
rect 576552 494292 576598 494448
rect 576810 495424 576856 495436
rect 576810 494448 576816 495424
rect 576850 494448 576856 495424
rect 576810 494436 576856 494448
rect 577068 495424 577114 495436
rect 577068 494448 577074 495424
rect 577108 494448 577114 495424
rect 576650 494398 576758 494404
rect 576650 494364 576662 494398
rect 576746 494364 576758 494398
rect 576650 494358 576758 494364
rect 576908 494398 577016 494404
rect 576908 494364 576920 494398
rect 577004 494364 577016 494398
rect 576908 494358 577016 494364
rect 577068 494292 577114 494448
rect 577326 495424 577372 495436
rect 577326 494448 577332 495424
rect 577366 494448 577372 495424
rect 577326 494436 577372 494448
rect 577584 495424 577630 495436
rect 577584 494448 577590 495424
rect 577624 494448 577630 495424
rect 577166 494398 577274 494404
rect 577166 494364 577178 494398
rect 577262 494364 577274 494398
rect 577166 494358 577274 494364
rect 577424 494398 577532 494404
rect 577424 494364 577436 494398
rect 577520 494364 577532 494398
rect 577424 494358 577532 494364
rect 577584 494292 577630 494448
rect 577698 495392 577744 495474
rect 577698 494418 577704 495392
rect 577738 494418 577744 495392
rect 577698 494406 577744 494418
rect 562120 494221 567614 494277
rect 562120 494161 562222 494221
rect 562282 494161 562342 494221
rect 562402 494161 562462 494221
rect 562522 494161 562582 494221
rect 562642 494161 562702 494221
rect 562762 494161 562822 494221
rect 562882 494161 562942 494221
rect 563002 494161 563062 494221
rect 563122 494161 563182 494221
rect 563242 494161 563302 494221
rect 563362 494161 563422 494221
rect 563482 494161 563542 494221
rect 563602 494161 563662 494221
rect 563722 494161 563782 494221
rect 563842 494161 563902 494221
rect 563962 494161 564022 494221
rect 564082 494161 564142 494221
rect 564202 494161 564262 494221
rect 564322 494161 564382 494221
rect 564442 494161 564502 494221
rect 564562 494161 564622 494221
rect 564682 494161 564742 494221
rect 564802 494161 564862 494221
rect 564922 494161 564982 494221
rect 565042 494161 565102 494221
rect 565162 494161 565222 494221
rect 565282 494161 565342 494221
rect 565402 494161 565462 494221
rect 565522 494161 565582 494221
rect 565642 494161 565702 494221
rect 565762 494161 565822 494221
rect 565882 494161 565942 494221
rect 566002 494161 566062 494221
rect 566122 494161 566182 494221
rect 566242 494161 566302 494221
rect 566362 494161 566422 494221
rect 566482 494161 566542 494221
rect 566602 494161 566662 494221
rect 566722 494161 566782 494221
rect 566842 494161 566902 494221
rect 566962 494161 567022 494221
rect 567082 494161 567142 494221
rect 567202 494161 567262 494221
rect 567322 494161 567382 494221
rect 567442 494161 567502 494221
rect 567562 494161 567614 494221
rect 562120 494101 567614 494161
rect 562120 494041 562222 494101
rect 562282 494041 562342 494101
rect 562402 494041 562462 494101
rect 562522 494041 562582 494101
rect 562642 494041 562702 494101
rect 562762 494041 562822 494101
rect 562882 494041 562942 494101
rect 563002 494041 563062 494101
rect 563122 494041 563182 494101
rect 563242 494041 563302 494101
rect 563362 494041 563422 494101
rect 563482 494041 563542 494101
rect 563602 494041 563662 494101
rect 563722 494041 563782 494101
rect 563842 494041 563902 494101
rect 563962 494041 564022 494101
rect 564082 494041 564142 494101
rect 564202 494041 564262 494101
rect 564322 494041 564382 494101
rect 564442 494041 564502 494101
rect 564562 494041 564622 494101
rect 564682 494041 564742 494101
rect 564802 494041 564862 494101
rect 564922 494041 564982 494101
rect 565042 494041 565102 494101
rect 565162 494041 565222 494101
rect 565282 494041 565342 494101
rect 565402 494041 565462 494101
rect 565522 494041 565582 494101
rect 565642 494041 565702 494101
rect 565762 494041 565822 494101
rect 565882 494041 565942 494101
rect 566002 494041 566062 494101
rect 566122 494041 566182 494101
rect 566242 494041 566302 494101
rect 566362 494041 566422 494101
rect 566482 494041 566542 494101
rect 566602 494041 566662 494101
rect 566722 494041 566782 494101
rect 566842 494041 566902 494101
rect 566962 494041 567022 494101
rect 567082 494041 567142 494101
rect 567202 494041 567262 494101
rect 567322 494041 567382 494101
rect 567442 494041 567502 494101
rect 567562 494041 567614 494101
rect 562120 494002 567614 494041
rect 572280 494236 577774 494292
rect 572280 494176 572332 494236
rect 572392 494176 572452 494236
rect 572512 494176 572572 494236
rect 572632 494176 572692 494236
rect 572752 494176 572812 494236
rect 572872 494176 572932 494236
rect 572992 494176 573052 494236
rect 573112 494176 573172 494236
rect 573232 494176 573292 494236
rect 573352 494176 573412 494236
rect 573472 494176 573532 494236
rect 573592 494176 573652 494236
rect 573712 494176 573772 494236
rect 573832 494176 573892 494236
rect 573952 494176 574012 494236
rect 574072 494176 574132 494236
rect 574192 494176 574252 494236
rect 574312 494176 574372 494236
rect 574432 494176 574492 494236
rect 574552 494176 574612 494236
rect 574672 494176 574732 494236
rect 574792 494176 574852 494236
rect 574912 494176 574972 494236
rect 575032 494176 575092 494236
rect 575152 494176 575212 494236
rect 575272 494176 575332 494236
rect 575392 494176 575452 494236
rect 575512 494176 575572 494236
rect 575632 494176 575692 494236
rect 575752 494176 575812 494236
rect 575872 494176 575932 494236
rect 575992 494176 576052 494236
rect 576112 494176 576172 494236
rect 576232 494176 576292 494236
rect 576352 494176 576412 494236
rect 576472 494176 576532 494236
rect 576592 494176 576652 494236
rect 576712 494176 576772 494236
rect 576832 494176 576892 494236
rect 576952 494176 577012 494236
rect 577072 494176 577132 494236
rect 577192 494176 577252 494236
rect 577312 494176 577372 494236
rect 577432 494176 577492 494236
rect 577552 494176 577612 494236
rect 577672 494176 577774 494236
rect 572280 494116 577774 494176
rect 572280 494056 572332 494116
rect 572392 494056 572452 494116
rect 572512 494056 572572 494116
rect 572632 494056 572692 494116
rect 572752 494056 572812 494116
rect 572872 494056 572932 494116
rect 572992 494056 573052 494116
rect 573112 494056 573172 494116
rect 573232 494056 573292 494116
rect 573352 494056 573412 494116
rect 573472 494056 573532 494116
rect 573592 494056 573652 494116
rect 573712 494056 573772 494116
rect 573832 494056 573892 494116
rect 573952 494056 574012 494116
rect 574072 494056 574132 494116
rect 574192 494056 574252 494116
rect 574312 494056 574372 494116
rect 574432 494056 574492 494116
rect 574552 494056 574612 494116
rect 574672 494056 574732 494116
rect 574792 494056 574852 494116
rect 574912 494056 574972 494116
rect 575032 494056 575092 494116
rect 575152 494056 575212 494116
rect 575272 494056 575332 494116
rect 575392 494056 575452 494116
rect 575512 494056 575572 494116
rect 575632 494056 575692 494116
rect 575752 494056 575812 494116
rect 575872 494056 575932 494116
rect 575992 494056 576052 494116
rect 576112 494056 576172 494116
rect 576232 494056 576292 494116
rect 576352 494056 576412 494116
rect 576472 494056 576532 494116
rect 576592 494056 576652 494116
rect 576712 494056 576772 494116
rect 576832 494056 576892 494116
rect 576952 494056 577012 494116
rect 577072 494056 577132 494116
rect 577192 494056 577252 494116
rect 577312 494056 577372 494116
rect 577432 494056 577492 494116
rect 577552 494056 577612 494116
rect 577672 494056 577774 494116
rect 572280 494017 577774 494056
rect 503900 475306 510526 475336
rect 503900 475206 503920 475306
rect 504020 475206 504144 475306
rect 504244 475206 504368 475306
rect 504468 475206 504592 475306
rect 504692 475206 504816 475306
rect 504916 475206 505040 475306
rect 505140 475206 505264 475306
rect 505364 475206 505488 475306
rect 505588 475206 505712 475306
rect 505812 475206 505936 475306
rect 506036 475206 506160 475306
rect 506260 475206 506384 475306
rect 506484 475206 506608 475306
rect 506708 475206 506832 475306
rect 506932 475206 507056 475306
rect 507156 475206 507280 475306
rect 507380 475206 507504 475306
rect 507604 475206 507728 475306
rect 507828 475206 507952 475306
rect 508052 475206 508176 475306
rect 508276 475206 508400 475306
rect 508500 475206 508624 475306
rect 508724 475206 508848 475306
rect 508948 475206 509072 475306
rect 509172 475206 509296 475306
rect 509396 475206 509520 475306
rect 509620 475206 509744 475306
rect 509844 475206 509968 475306
rect 510068 475206 510192 475306
rect 510292 475206 510416 475306
rect 510516 475206 510526 475306
rect 503900 475082 510526 475206
rect 503900 474982 503920 475082
rect 504020 474982 504144 475082
rect 504244 474982 504368 475082
rect 504468 474982 504592 475082
rect 504692 474982 504816 475082
rect 504916 474982 505040 475082
rect 505140 474982 505264 475082
rect 505364 474982 505488 475082
rect 505588 474982 505712 475082
rect 505812 474982 505936 475082
rect 506036 474982 506160 475082
rect 506260 474982 506384 475082
rect 506484 474982 506608 475082
rect 506708 474982 506832 475082
rect 506932 474982 507056 475082
rect 507156 474982 507280 475082
rect 507380 474982 507504 475082
rect 507604 474982 507728 475082
rect 507828 474982 507952 475082
rect 508052 474982 508176 475082
rect 508276 474982 508400 475082
rect 508500 474982 508624 475082
rect 508724 474982 508848 475082
rect 508948 474982 509072 475082
rect 509172 474982 509296 475082
rect 509396 474982 509520 475082
rect 509620 474982 509744 475082
rect 509844 474982 509968 475082
rect 510068 474982 510192 475082
rect 510292 474982 510416 475082
rect 510516 474982 510526 475082
rect 503900 474858 510526 474982
rect 503900 474758 503920 474858
rect 504020 474758 504144 474858
rect 504244 474758 504368 474858
rect 504468 474758 504592 474858
rect 504692 474758 504816 474858
rect 504916 474758 505040 474858
rect 505140 474758 505264 474858
rect 505364 474758 505488 474858
rect 505588 474758 505712 474858
rect 505812 474758 505936 474858
rect 506036 474758 506160 474858
rect 506260 474758 506384 474858
rect 506484 474758 506608 474858
rect 506708 474758 506832 474858
rect 506932 474758 507056 474858
rect 507156 474758 507280 474858
rect 507380 474758 507504 474858
rect 507604 474758 507728 474858
rect 507828 474758 507952 474858
rect 508052 474758 508176 474858
rect 508276 474758 508400 474858
rect 508500 474758 508624 474858
rect 508724 474758 508848 474858
rect 508948 474758 509072 474858
rect 509172 474758 509296 474858
rect 509396 474758 509520 474858
rect 509620 474758 509744 474858
rect 509844 474758 509968 474858
rect 510068 474758 510192 474858
rect 510292 474758 510416 474858
rect 510516 474758 510526 474858
rect 503900 474634 510526 474758
rect 503900 474534 503920 474634
rect 504020 474534 504144 474634
rect 504244 474534 504368 474634
rect 504468 474534 504592 474634
rect 504692 474534 504816 474634
rect 504916 474534 505040 474634
rect 505140 474534 505264 474634
rect 505364 474534 505488 474634
rect 505588 474534 505712 474634
rect 505812 474534 505936 474634
rect 506036 474534 506160 474634
rect 506260 474534 506384 474634
rect 506484 474534 506608 474634
rect 506708 474534 506832 474634
rect 506932 474534 507056 474634
rect 507156 474534 507280 474634
rect 507380 474534 507504 474634
rect 507604 474534 507728 474634
rect 507828 474534 507952 474634
rect 508052 474534 508176 474634
rect 508276 474534 508400 474634
rect 508500 474534 508624 474634
rect 508724 474534 508848 474634
rect 508948 474534 509072 474634
rect 509172 474534 509296 474634
rect 509396 474534 509520 474634
rect 509620 474534 509744 474634
rect 509844 474534 509968 474634
rect 510068 474534 510192 474634
rect 510292 474534 510416 474634
rect 510516 474534 510526 474634
rect 503900 474410 510526 474534
rect 500364 474280 501424 474320
rect 500364 474180 500398 474280
rect 500498 474180 500622 474280
rect 500722 474180 500846 474280
rect 500946 474180 501070 474280
rect 501170 474180 501294 474280
rect 501394 474180 501424 474280
rect 503900 474310 503920 474410
rect 504020 474310 504144 474410
rect 504244 474310 504368 474410
rect 504468 474310 504592 474410
rect 504692 474310 504816 474410
rect 504916 474310 505040 474410
rect 505140 474310 505264 474410
rect 505364 474310 505488 474410
rect 505588 474310 505712 474410
rect 505812 474310 505936 474410
rect 506036 474310 506160 474410
rect 506260 474310 506384 474410
rect 506484 474310 506608 474410
rect 506708 474310 506832 474410
rect 506932 474310 507056 474410
rect 507156 474310 507280 474410
rect 507380 474310 507504 474410
rect 507604 474310 507728 474410
rect 507828 474310 507952 474410
rect 508052 474310 508176 474410
rect 508276 474310 508400 474410
rect 508500 474310 508624 474410
rect 508724 474310 508848 474410
rect 508948 474310 509072 474410
rect 509172 474310 509296 474410
rect 509396 474310 509520 474410
rect 509620 474310 509744 474410
rect 509844 474310 509968 474410
rect 510068 474310 510192 474410
rect 510292 474310 510416 474410
rect 510516 474310 510526 474410
rect 503900 474278 510526 474310
rect 517280 475306 523940 475336
rect 517280 475206 517320 475306
rect 517420 475206 517544 475306
rect 517644 475206 517768 475306
rect 517868 475206 517992 475306
rect 518092 475206 518216 475306
rect 518316 475206 518440 475306
rect 518540 475206 518664 475306
rect 518764 475206 518888 475306
rect 518988 475206 519112 475306
rect 519212 475206 519336 475306
rect 519436 475206 519560 475306
rect 519660 475206 519784 475306
rect 519884 475206 520008 475306
rect 520108 475206 520232 475306
rect 520332 475206 520456 475306
rect 520556 475206 520680 475306
rect 520780 475206 520904 475306
rect 521004 475206 521128 475306
rect 521228 475206 521352 475306
rect 521452 475206 521576 475306
rect 521676 475206 521800 475306
rect 521900 475206 522024 475306
rect 522124 475206 522248 475306
rect 522348 475206 522472 475306
rect 522572 475206 522696 475306
rect 522796 475206 522920 475306
rect 523020 475206 523144 475306
rect 523244 475206 523368 475306
rect 523468 475206 523592 475306
rect 523692 475206 523816 475306
rect 523916 475206 523940 475306
rect 517280 475082 523940 475206
rect 517280 474982 517320 475082
rect 517420 474982 517544 475082
rect 517644 474982 517768 475082
rect 517868 474982 517992 475082
rect 518092 474982 518216 475082
rect 518316 474982 518440 475082
rect 518540 474982 518664 475082
rect 518764 474982 518888 475082
rect 518988 474982 519112 475082
rect 519212 474982 519336 475082
rect 519436 474982 519560 475082
rect 519660 474982 519784 475082
rect 519884 474982 520008 475082
rect 520108 474982 520232 475082
rect 520332 474982 520456 475082
rect 520556 474982 520680 475082
rect 520780 474982 520904 475082
rect 521004 474982 521128 475082
rect 521228 474982 521352 475082
rect 521452 474982 521576 475082
rect 521676 474982 521800 475082
rect 521900 474982 522024 475082
rect 522124 474982 522248 475082
rect 522348 474982 522472 475082
rect 522572 474982 522696 475082
rect 522796 474982 522920 475082
rect 523020 474982 523144 475082
rect 523244 474982 523368 475082
rect 523468 474982 523592 475082
rect 523692 474982 523816 475082
rect 523916 474982 523940 475082
rect 517280 474858 523940 474982
rect 517280 474758 517320 474858
rect 517420 474758 517544 474858
rect 517644 474758 517768 474858
rect 517868 474758 517992 474858
rect 518092 474758 518216 474858
rect 518316 474758 518440 474858
rect 518540 474758 518664 474858
rect 518764 474758 518888 474858
rect 518988 474758 519112 474858
rect 519212 474758 519336 474858
rect 519436 474758 519560 474858
rect 519660 474758 519784 474858
rect 519884 474758 520008 474858
rect 520108 474758 520232 474858
rect 520332 474758 520456 474858
rect 520556 474758 520680 474858
rect 520780 474758 520904 474858
rect 521004 474758 521128 474858
rect 521228 474758 521352 474858
rect 521452 474758 521576 474858
rect 521676 474758 521800 474858
rect 521900 474758 522024 474858
rect 522124 474758 522248 474858
rect 522348 474758 522472 474858
rect 522572 474758 522696 474858
rect 522796 474758 522920 474858
rect 523020 474758 523144 474858
rect 523244 474758 523368 474858
rect 523468 474758 523592 474858
rect 523692 474758 523816 474858
rect 523916 474758 523940 474858
rect 517280 474634 523940 474758
rect 517280 474534 517320 474634
rect 517420 474534 517544 474634
rect 517644 474534 517768 474634
rect 517868 474534 517992 474634
rect 518092 474534 518216 474634
rect 518316 474534 518440 474634
rect 518540 474534 518664 474634
rect 518764 474534 518888 474634
rect 518988 474534 519112 474634
rect 519212 474534 519336 474634
rect 519436 474534 519560 474634
rect 519660 474534 519784 474634
rect 519884 474534 520008 474634
rect 520108 474534 520232 474634
rect 520332 474534 520456 474634
rect 520556 474534 520680 474634
rect 520780 474534 520904 474634
rect 521004 474534 521128 474634
rect 521228 474534 521352 474634
rect 521452 474534 521576 474634
rect 521676 474534 521800 474634
rect 521900 474534 522024 474634
rect 522124 474534 522248 474634
rect 522348 474534 522472 474634
rect 522572 474534 522696 474634
rect 522796 474534 522920 474634
rect 523020 474534 523144 474634
rect 523244 474534 523368 474634
rect 523468 474534 523592 474634
rect 523692 474534 523816 474634
rect 523916 474534 523940 474634
rect 517280 474410 523940 474534
rect 517280 474310 517320 474410
rect 517420 474310 517544 474410
rect 517644 474310 517768 474410
rect 517868 474310 517992 474410
rect 518092 474310 518216 474410
rect 518316 474310 518440 474410
rect 518540 474310 518664 474410
rect 518764 474310 518888 474410
rect 518988 474310 519112 474410
rect 519212 474310 519336 474410
rect 519436 474310 519560 474410
rect 519660 474310 519784 474410
rect 519884 474310 520008 474410
rect 520108 474310 520232 474410
rect 520332 474310 520456 474410
rect 520556 474310 520680 474410
rect 520780 474310 520904 474410
rect 521004 474310 521128 474410
rect 521228 474310 521352 474410
rect 521452 474310 521576 474410
rect 521676 474310 521800 474410
rect 521900 474310 522024 474410
rect 522124 474310 522248 474410
rect 522348 474310 522472 474410
rect 522572 474310 522696 474410
rect 522796 474310 522920 474410
rect 523020 474310 523144 474410
rect 523244 474310 523368 474410
rect 523468 474310 523592 474410
rect 523692 474310 523816 474410
rect 523916 474310 523940 474410
rect 517280 474276 523940 474310
rect 527584 474280 528644 474320
rect 500364 474056 501424 474180
rect 500364 473956 500398 474056
rect 500498 473956 500622 474056
rect 500722 473956 500846 474056
rect 500946 473956 501070 474056
rect 501170 473956 501294 474056
rect 501394 473956 501424 474056
rect 500364 473832 501424 473956
rect 500364 473732 500398 473832
rect 500498 473732 500622 473832
rect 500722 473732 500846 473832
rect 500946 473732 501070 473832
rect 501170 473732 501294 473832
rect 501394 473732 501424 473832
rect 500364 473608 501424 473732
rect 500364 473508 500398 473608
rect 500498 473508 500622 473608
rect 500722 473508 500846 473608
rect 500946 473508 501070 473608
rect 501170 473508 501294 473608
rect 501394 473508 501424 473608
rect 500364 473384 501424 473508
rect 500364 473284 500398 473384
rect 500498 473284 500622 473384
rect 500722 473284 500846 473384
rect 500946 473284 501070 473384
rect 501170 473284 501294 473384
rect 501394 473284 501424 473384
rect 500364 473160 501424 473284
rect 500364 473060 500398 473160
rect 500498 473060 500622 473160
rect 500722 473060 500846 473160
rect 500946 473060 501070 473160
rect 501170 473060 501294 473160
rect 501394 473060 501424 473160
rect 500364 472936 501424 473060
rect 500364 472836 500398 472936
rect 500498 472836 500622 472936
rect 500722 472836 500846 472936
rect 500946 472836 501070 472936
rect 501170 472836 501294 472936
rect 501394 472836 501424 472936
rect 500364 472712 501424 472836
rect 527584 474180 527618 474280
rect 527718 474180 527842 474280
rect 527942 474180 528066 474280
rect 528166 474180 528290 474280
rect 528390 474180 528514 474280
rect 528614 474180 528644 474280
rect 527584 474056 528644 474180
rect 527584 473956 527618 474056
rect 527718 473956 527842 474056
rect 527942 473956 528066 474056
rect 528166 473956 528290 474056
rect 528390 473956 528514 474056
rect 528614 473956 528644 474056
rect 527584 473832 528644 473956
rect 527584 473732 527618 473832
rect 527718 473732 527842 473832
rect 527942 473732 528066 473832
rect 528166 473732 528290 473832
rect 528390 473732 528514 473832
rect 528614 473732 528644 473832
rect 527584 473608 528644 473732
rect 527584 473508 527618 473608
rect 527718 473508 527842 473608
rect 527942 473508 528066 473608
rect 528166 473508 528290 473608
rect 528390 473508 528514 473608
rect 528614 473508 528644 473608
rect 527584 473384 528644 473508
rect 527584 473284 527618 473384
rect 527718 473284 527842 473384
rect 527942 473284 528066 473384
rect 528166 473284 528290 473384
rect 528390 473284 528514 473384
rect 528614 473284 528644 473384
rect 527584 473160 528644 473284
rect 527584 473060 527618 473160
rect 527718 473060 527842 473160
rect 527942 473060 528066 473160
rect 528166 473060 528290 473160
rect 528390 473060 528514 473160
rect 528614 473060 528644 473160
rect 527584 472936 528644 473060
rect 527584 472836 527618 472936
rect 527718 472836 527842 472936
rect 527942 472836 528066 472936
rect 528166 472836 528290 472936
rect 528390 472836 528514 472936
rect 528614 472836 528644 472936
rect 506558 472764 506958 472770
rect 506558 472730 506570 472764
rect 506946 472730 506958 472764
rect 506558 472724 506958 472730
rect 500364 472612 500398 472712
rect 500498 472612 500622 472712
rect 500722 472612 500846 472712
rect 500946 472612 501070 472712
rect 501170 472612 501294 472712
rect 501394 472612 501424 472712
rect 527584 472712 528644 472836
rect 500364 472488 501424 472612
rect 500364 472388 500398 472488
rect 500498 472388 500622 472488
rect 500722 472388 500846 472488
rect 500946 472388 501070 472488
rect 501170 472388 501294 472488
rect 501394 472388 501424 472488
rect 506990 472610 507036 472622
rect 506990 472426 506996 472610
rect 507030 472426 507036 472610
rect 527584 472612 527618 472712
rect 527718 472612 527842 472712
rect 527942 472612 528066 472712
rect 528166 472612 528290 472712
rect 528390 472612 528514 472712
rect 528614 472612 528644 472712
rect 506990 472414 507036 472426
rect 525660 472498 526498 472504
rect 500364 472264 501424 472388
rect 500364 472164 500398 472264
rect 500498 472164 500622 472264
rect 500722 472164 500846 472264
rect 500946 472164 501070 472264
rect 501170 472164 501294 472264
rect 501394 472164 501424 472264
rect 506364 472316 506428 472322
rect 506364 472264 506370 472316
rect 506422 472312 506428 472316
rect 506422 472306 507030 472312
rect 506422 472272 506570 472306
rect 506946 472272 507030 472306
rect 506422 472268 507030 472272
rect 506422 472266 506958 472268
rect 506422 472264 506428 472266
rect 506364 472258 506428 472264
rect 506996 472176 507030 472268
rect 500364 472040 501424 472164
rect 500364 471940 500398 472040
rect 500498 471940 500622 472040
rect 500722 471940 500846 472040
rect 500946 471940 501070 472040
rect 501170 471940 501294 472040
rect 501394 471940 501424 472040
rect 506978 472152 507042 472176
rect 506978 471968 506996 472152
rect 507030 471968 507042 472152
rect 506978 471944 507042 471968
rect 500364 471816 501424 471940
rect 507082 471858 507158 471870
rect 507082 471854 507094 471858
rect 500364 471716 500398 471816
rect 500498 471716 500622 471816
rect 500722 471716 500846 471816
rect 500946 471716 501070 471816
rect 501170 471716 501294 471816
rect 501394 471716 501424 471816
rect 506558 471848 507094 471854
rect 506558 471814 506570 471848
rect 506946 471814 507094 471848
rect 506558 471808 507094 471814
rect 507082 471806 507094 471808
rect 507146 471806 507158 471858
rect 507082 471794 507158 471806
rect 500364 471592 501424 471716
rect 500364 471492 500398 471592
rect 500498 471492 500622 471592
rect 500722 471492 500846 471592
rect 500946 471492 501070 471592
rect 501170 471492 501294 471592
rect 501394 471492 501424 471592
rect 506990 471694 507036 471706
rect 506990 471510 506996 471694
rect 507030 471510 507036 471694
rect 506990 471498 507036 471510
rect 500364 471368 501424 471492
rect 500364 471268 500398 471368
rect 500498 471268 500622 471368
rect 500722 471268 500846 471368
rect 500946 471268 501070 471368
rect 501170 471268 501294 471368
rect 501394 471268 501424 471368
rect 506158 471398 506222 471404
rect 506158 471346 506164 471398
rect 506216 471396 506222 471398
rect 506216 471390 506958 471396
rect 506216 471356 506570 471390
rect 506946 471356 506958 471390
rect 506216 471350 506958 471356
rect 506216 471346 506222 471350
rect 506158 471340 506222 471346
rect 500364 471144 501424 471268
rect 500364 471044 500398 471144
rect 500498 471044 500622 471144
rect 500722 471044 500846 471144
rect 500946 471044 501070 471144
rect 501170 471044 501294 471144
rect 501394 471044 501424 471144
rect 500364 470920 501424 471044
rect 506990 471236 507036 471248
rect 506990 471052 506996 471236
rect 507030 471052 507036 471236
rect 506990 471040 507036 471052
rect 507082 470942 507158 470954
rect 507082 470938 507094 470942
rect 500364 470820 500398 470920
rect 500498 470820 500622 470920
rect 500722 470820 500846 470920
rect 500946 470820 501070 470920
rect 501170 470820 501294 470920
rect 501394 470820 501424 470920
rect 506558 470932 507094 470938
rect 506558 470898 506570 470932
rect 506946 470898 507094 470932
rect 506558 470892 507094 470898
rect 507082 470890 507094 470892
rect 507146 470890 507158 470942
rect 507082 470878 507158 470890
rect 500364 470696 501424 470820
rect 500364 470596 500398 470696
rect 500498 470596 500622 470696
rect 500722 470596 500846 470696
rect 500946 470596 501070 470696
rect 501170 470596 501294 470696
rect 501394 470596 501424 470696
rect 500364 470472 501424 470596
rect 506978 470778 507042 470812
rect 506978 470594 506996 470778
rect 507030 470594 507042 470778
rect 506978 470580 507042 470594
rect 500364 470372 500398 470472
rect 500498 470372 500622 470472
rect 500722 470372 500846 470472
rect 500946 470372 501070 470472
rect 501170 470372 501294 470472
rect 501394 470372 501424 470472
rect 506370 470482 506434 470488
rect 506370 470430 506376 470482
rect 506428 470480 506434 470482
rect 506996 470480 507030 470580
rect 506428 470474 507030 470480
rect 506428 470440 506570 470474
rect 506946 470440 507030 470474
rect 506428 470434 507030 470440
rect 506428 470430 506434 470434
rect 506370 470424 506434 470430
rect 500364 470248 501424 470372
rect 500364 470148 500398 470248
rect 500498 470148 500622 470248
rect 500722 470148 500846 470248
rect 500946 470148 501070 470248
rect 501170 470148 501294 470248
rect 501394 470148 501424 470248
rect 506990 470320 507036 470332
rect 500364 470024 501424 470148
rect 502864 470202 505580 470218
rect 502864 470192 503226 470202
rect 502864 470140 502874 470192
rect 502978 470140 503226 470192
rect 502864 470102 503226 470140
rect 505568 470102 505580 470202
rect 506990 470136 506996 470320
rect 507030 470136 507036 470320
rect 506990 470124 507036 470136
rect 509928 470184 510136 470206
rect 509928 470124 509940 470184
rect 510010 470124 510034 470184
rect 510104 470124 510136 470184
rect 502864 470086 505580 470102
rect 509928 470112 510136 470124
rect 500364 469924 500398 470024
rect 500498 469924 500622 470024
rect 500722 469924 500846 470024
rect 500946 469924 501070 470024
rect 501170 469924 501294 470024
rect 501394 469924 501424 470024
rect 509928 470052 509940 470112
rect 510010 470052 510034 470112
rect 510104 470052 510136 470112
rect 509928 470040 510136 470052
rect 506558 470016 506958 470022
rect 506558 469982 506570 470016
rect 506946 469982 506958 470016
rect 506558 469976 506958 469982
rect 509928 469980 509940 470040
rect 510010 469980 510034 470040
rect 510104 469980 510136 470040
rect 500364 469800 501424 469924
rect 509928 469968 510136 469980
rect 509928 469908 509940 469968
rect 510010 469908 510034 469968
rect 510104 469908 510136 469968
rect 509928 469896 510136 469908
rect 500364 469700 500398 469800
rect 500498 469700 500622 469800
rect 500722 469700 500846 469800
rect 500946 469700 501070 469800
rect 501170 469700 501294 469800
rect 501394 469700 501424 469800
rect 500364 469576 501424 469700
rect 502664 469876 506434 469882
rect 502664 469682 502670 469876
rect 502784 469682 506370 469876
rect 506428 469682 506434 469876
rect 502664 469676 506434 469682
rect 509928 469836 509940 469896
rect 510010 469836 510034 469896
rect 510104 469836 510136 469896
rect 509928 469824 510136 469836
rect 509928 469764 509940 469824
rect 510010 469764 510034 469824
rect 510104 469764 510136 469824
rect 509928 469752 510136 469764
rect 509928 469692 509940 469752
rect 510010 469692 510034 469752
rect 510104 469692 510136 469752
rect 509928 469680 510136 469692
rect 509928 469620 509940 469680
rect 510010 469620 510034 469680
rect 510104 469620 510136 469680
rect 500364 469476 500398 469576
rect 500498 469476 500622 469576
rect 500722 469476 500846 469576
rect 500946 469476 501070 469576
rect 501170 469476 501294 469576
rect 501394 469476 501424 469576
rect 502864 469570 502988 469580
rect 502864 469518 502874 469570
rect 502978 469566 502988 469570
rect 502978 469560 505756 469566
rect 502978 469526 503100 469560
rect 505656 469526 505756 469560
rect 502978 469520 505756 469526
rect 502978 469518 502988 469520
rect 502864 469508 502988 469518
rect 500364 469352 501424 469476
rect 500364 469252 500398 469352
rect 500498 469252 500622 469352
rect 500722 469252 500846 469352
rect 500946 469252 501070 469352
rect 501170 469252 501294 469352
rect 501394 469252 501424 469352
rect 500364 469128 501424 469252
rect 500364 469028 500398 469128
rect 500498 469028 500622 469128
rect 500722 469028 500846 469128
rect 500946 469028 501070 469128
rect 501170 469028 501294 469128
rect 501394 469028 501424 469128
rect 505708 469406 505756 469520
rect 505708 469222 505715 469406
rect 505749 469222 505756 469406
rect 502864 469112 502988 469122
rect 502864 469060 502874 469112
rect 502978 469108 502988 469112
rect 505708 469108 505756 469222
rect 502978 469102 505756 469108
rect 502978 469068 503100 469102
rect 505656 469068 505756 469102
rect 502978 469062 505756 469068
rect 502978 469060 502988 469062
rect 502864 469050 502988 469060
rect 500364 468904 501424 469028
rect 502664 468996 502788 469006
rect 502664 468944 502674 468996
rect 502778 468992 502788 468996
rect 503088 468992 505668 468994
rect 502778 468988 505668 468992
rect 502778 468954 503100 468988
rect 505656 468954 505668 468988
rect 502778 468950 505668 468954
rect 502778 468944 502788 468950
rect 503088 468948 505668 468950
rect 502664 468934 502788 468944
rect 500364 468804 500398 468904
rect 500498 468804 500622 468904
rect 500722 468804 500846 468904
rect 500946 468804 501070 468904
rect 501170 468804 501294 468904
rect 501394 468804 501424 468904
rect 500364 468680 501424 468804
rect 500364 468580 500398 468680
rect 500498 468580 500622 468680
rect 500722 468580 500846 468680
rect 500946 468580 501070 468680
rect 501170 468580 501294 468680
rect 501394 468580 501424 468680
rect 505708 468834 509820 468846
rect 505708 468650 505715 468834
rect 505749 468720 509820 468834
rect 505749 468668 505802 468720
rect 506056 468668 509820 468720
rect 505749 468650 509820 468668
rect 505708 468638 509820 468650
rect 500364 468456 501424 468580
rect 502864 468536 502988 468546
rect 502864 468484 502874 468536
rect 502978 468530 502988 468536
rect 503088 468530 505668 468536
rect 502978 468496 503100 468530
rect 505656 468496 505668 468530
rect 502978 468484 502988 468496
rect 503088 468490 505668 468496
rect 502864 468474 502988 468484
rect 500364 468356 500398 468456
rect 500498 468356 500622 468456
rect 500722 468356 500846 468456
rect 500946 468356 501070 468456
rect 501170 468356 501294 468456
rect 501394 468356 501424 468456
rect 502664 468424 502788 468434
rect 502664 468372 502674 468424
rect 502778 468420 502788 468424
rect 503088 468420 505668 468422
rect 502778 468416 505668 468420
rect 502778 468382 503100 468416
rect 505656 468382 505668 468416
rect 502778 468378 505668 468382
rect 502778 468372 502788 468378
rect 503088 468376 505668 468378
rect 506452 468392 508084 468402
rect 506452 468386 508158 468392
rect 502664 468362 502788 468372
rect 500364 468232 501424 468356
rect 506452 468286 506470 468386
rect 508068 468286 508158 468386
rect 500364 468132 500398 468232
rect 500498 468132 500622 468232
rect 500722 468132 500846 468232
rect 500946 468132 501070 468232
rect 501170 468132 501294 468232
rect 501394 468132 501424 468232
rect 500364 468008 501424 468132
rect 505708 468262 506062 468286
rect 506452 468278 508158 468286
rect 506452 468270 508084 468278
rect 505708 468078 505715 468262
rect 505749 468160 506062 468262
rect 505749 468108 505802 468160
rect 506056 468108 506062 468160
rect 505749 468078 506062 468108
rect 505709 468066 505755 468078
rect 500364 467908 500398 468008
rect 500498 467908 500622 468008
rect 500722 467908 500846 468008
rect 500946 467908 501070 468008
rect 501170 467908 501294 468008
rect 501394 467908 501424 468008
rect 500364 467784 501424 467908
rect 502864 467964 502988 467974
rect 502864 467912 502874 467964
rect 502978 467958 502988 467964
rect 503088 467958 505668 467964
rect 502978 467924 503100 467958
rect 505656 467924 505668 467958
rect 502978 467918 505668 467924
rect 502978 467916 505652 467918
rect 502978 467912 502988 467916
rect 502864 467902 502988 467912
rect 502664 467852 502788 467862
rect 502664 467800 502674 467852
rect 502778 467848 502788 467852
rect 503088 467848 505668 467850
rect 502778 467844 505668 467848
rect 502778 467810 503100 467844
rect 505656 467810 505668 467844
rect 508112 467840 508158 468278
rect 502778 467806 505668 467810
rect 502778 467800 502788 467806
rect 503088 467804 505668 467806
rect 506280 467834 508158 467840
rect 502664 467790 502788 467800
rect 506280 467800 506292 467834
rect 508068 467800 508158 467834
rect 506280 467794 508158 467800
rect 500364 467684 500398 467784
rect 500498 467684 500622 467784
rect 500722 467684 500846 467784
rect 500946 467684 501070 467784
rect 501170 467684 501294 467784
rect 501394 467684 501424 467784
rect 500364 467660 501424 467684
rect 505708 467690 506062 467726
rect 505708 467518 505715 467690
rect 505709 467506 505715 467518
rect 505749 467600 506062 467690
rect 505749 467548 505802 467600
rect 506056 467548 506062 467600
rect 505749 467518 506062 467548
rect 508112 467680 508158 467794
rect 505749 467506 505755 467518
rect 505709 467494 505755 467506
rect 508112 467496 508118 467680
rect 508152 467496 508158 467680
rect 502864 467392 502988 467402
rect 502864 467340 502874 467392
rect 502978 467386 502988 467392
rect 503088 467386 505668 467392
rect 502978 467352 503100 467386
rect 505656 467352 505668 467386
rect 508112 467382 508158 467496
rect 502978 467346 505668 467352
rect 506280 467376 508158 467382
rect 502978 467340 505652 467346
rect 502864 467336 505652 467340
rect 506280 467342 506292 467376
rect 508068 467342 508158 467376
rect 506280 467336 508158 467342
rect 509464 468128 509820 468638
rect 509928 468200 510136 469620
rect 509928 468166 509940 468200
rect 510124 468166 510136 468200
rect 509928 468160 510136 468166
rect 510258 468840 510826 468852
rect 510258 468128 510470 468840
rect 509464 468116 509826 468128
rect 502864 467330 502988 467336
rect 503088 467272 505668 467278
rect 503088 467238 503100 467272
rect 505656 467264 505668 467272
rect 506280 467264 508080 467268
rect 505656 467262 508080 467264
rect 505656 467238 506292 467262
rect 503088 467232 506292 467238
rect 505652 467230 506292 467232
rect 505710 467130 505750 467230
rect 506280 467228 506292 467230
rect 508068 467228 508080 467262
rect 506280 467222 508080 467228
rect 505709 467128 505755 467130
rect 505698 467122 505768 467128
rect 505698 466914 505708 467122
rect 505766 466914 505768 467122
rect 505698 466908 505768 466914
rect 508112 467108 508158 467120
rect 508112 466924 508118 467108
rect 508152 467088 508292 467108
rect 508152 466944 508218 467088
rect 508272 466944 508292 467088
rect 508152 466924 508292 466944
rect 508112 466912 508158 466924
rect 502864 466820 502988 466830
rect 502864 466768 502874 466820
rect 502978 466814 502988 466820
rect 503088 466814 505668 466820
rect 505710 466818 505746 466908
rect 506092 466820 506216 466830
rect 502978 466780 503100 466814
rect 505656 466780 505668 466814
rect 502978 466774 505668 466780
rect 502978 466772 505652 466774
rect 502978 466768 502988 466772
rect 502864 466758 502988 466768
rect 506092 466768 506102 466820
rect 506206 466804 506216 466820
rect 506280 466804 508080 466810
rect 506206 466770 506292 466804
rect 508068 466770 508080 466804
rect 506206 466768 506216 466770
rect 506092 466758 506216 466768
rect 506280 466764 508080 466770
rect 503088 466700 505668 466706
rect 503088 466666 503100 466700
rect 505656 466692 505668 466700
rect 505796 466700 506062 466706
rect 505796 466692 505802 466700
rect 505656 466666 505802 466692
rect 503088 466660 505802 466666
rect 505656 466658 505802 466660
rect 505796 466648 505802 466658
rect 506056 466692 506062 466700
rect 506280 466692 508080 466696
rect 506056 466690 508080 466692
rect 506056 466658 506292 466690
rect 506056 466648 506062 466658
rect 506280 466656 506292 466658
rect 508068 466656 508080 466690
rect 506280 466650 508080 466656
rect 505796 466642 506062 466648
rect 502606 466620 502738 466632
rect 502606 464278 502622 466620
rect 502722 464278 502738 466620
rect 505709 466556 505755 466558
rect 505698 466550 505768 466556
rect 505698 466342 505704 466550
rect 505762 466342 505768 466550
rect 505698 466336 505768 466342
rect 508112 466536 508158 466548
rect 508112 466352 508118 466536
rect 508152 466516 508432 466536
rect 508152 466372 508358 466516
rect 508412 466372 508432 466516
rect 508152 466352 508432 466372
rect 508112 466340 508158 466352
rect 502864 466248 502988 466258
rect 506092 466248 506216 466258
rect 502864 466196 502874 466248
rect 502978 466242 502988 466248
rect 503088 466242 505668 466248
rect 502978 466208 503100 466242
rect 505656 466208 505668 466242
rect 502978 466202 505668 466208
rect 502978 466200 505652 466202
rect 502978 466196 502988 466200
rect 502864 466186 502988 466196
rect 506092 466196 506102 466248
rect 506206 466232 506216 466248
rect 506280 466232 508080 466238
rect 506206 466198 506292 466232
rect 508068 466198 508080 466232
rect 506206 466196 506216 466198
rect 506092 466186 506216 466196
rect 506280 466192 508080 466198
rect 503088 466128 505668 466134
rect 503088 466094 503100 466128
rect 505656 466120 505668 466128
rect 506280 466120 508080 466124
rect 505656 466118 508080 466120
rect 505656 466094 506292 466118
rect 503088 466088 506292 466094
rect 505656 466086 506292 466088
rect 505714 465986 505750 466086
rect 506280 466084 506292 466086
rect 508068 466084 508080 466118
rect 506280 466078 508080 466084
rect 505709 465984 505755 465986
rect 505702 465978 505772 465984
rect 505702 465770 505708 465978
rect 505766 465770 505772 465978
rect 505702 465764 505772 465770
rect 508112 465964 508158 465976
rect 508112 465780 508118 465964
rect 508152 465944 508292 465964
rect 508152 465800 508218 465944
rect 508272 465800 508292 465944
rect 508152 465780 508292 465800
rect 508112 465768 508158 465780
rect 502864 465676 502988 465686
rect 502864 465624 502874 465676
rect 502978 465670 502988 465676
rect 503088 465670 505668 465676
rect 505714 465674 505750 465764
rect 506092 465676 506216 465686
rect 502978 465636 503100 465670
rect 505656 465636 505668 465670
rect 502978 465624 502988 465636
rect 503088 465630 505668 465636
rect 502864 465614 502988 465624
rect 506092 465624 506102 465676
rect 506206 465660 506216 465676
rect 506280 465660 508080 465666
rect 506206 465626 506292 465660
rect 508068 465626 508080 465660
rect 506206 465624 506216 465626
rect 506092 465614 506216 465624
rect 506280 465620 508080 465626
rect 503088 465556 505668 465562
rect 503088 465522 503100 465556
rect 505656 465548 505668 465556
rect 505796 465556 506062 465562
rect 505796 465548 505802 465556
rect 505656 465522 505802 465548
rect 503088 465516 505802 465522
rect 505656 465514 505802 465516
rect 505796 465504 505802 465514
rect 506056 465548 506062 465556
rect 506280 465548 508080 465552
rect 506056 465546 508080 465548
rect 506056 465514 506292 465546
rect 506056 465504 506062 465514
rect 506280 465512 506292 465514
rect 508068 465512 508080 465546
rect 506280 465506 508080 465512
rect 505796 465498 506062 465504
rect 505709 465412 505755 465414
rect 505702 465406 505772 465412
rect 505702 465198 505708 465406
rect 505766 465198 505772 465406
rect 505702 465192 505772 465198
rect 508112 465392 508158 465404
rect 508112 465208 508118 465392
rect 508152 465372 508432 465392
rect 508152 465228 508358 465372
rect 508412 465228 508432 465372
rect 508152 465208 508432 465228
rect 508112 465196 508158 465208
rect 502864 465104 502988 465114
rect 506092 465104 506216 465114
rect 502864 465052 502874 465104
rect 502978 465098 502988 465104
rect 503088 465098 505668 465104
rect 502978 465064 503100 465098
rect 505656 465064 505668 465098
rect 502978 465052 502988 465064
rect 503088 465058 505668 465064
rect 502864 465042 502988 465052
rect 506092 465052 506102 465104
rect 506206 465088 506216 465104
rect 506280 465088 508080 465094
rect 506206 465054 506292 465088
rect 508068 465054 508080 465088
rect 506206 465052 506216 465054
rect 506092 465042 506216 465052
rect 506280 465048 508080 465054
rect 503088 464984 505668 464990
rect 503088 464950 503100 464984
rect 505656 464976 505668 464984
rect 506280 464976 508080 464980
rect 505656 464974 508080 464976
rect 505656 464950 506292 464974
rect 503088 464944 506292 464950
rect 505656 464942 506292 464944
rect 505714 464842 505750 464942
rect 506280 464940 506292 464942
rect 508068 464940 508080 464974
rect 506280 464934 508080 464940
rect 505709 464840 505755 464842
rect 505702 464834 505772 464840
rect 505702 464626 505708 464834
rect 505766 464626 505772 464834
rect 505702 464620 505772 464626
rect 508112 464820 508158 464832
rect 508112 464636 508118 464820
rect 508152 464800 508292 464820
rect 508152 464656 508218 464800
rect 508272 464656 508292 464800
rect 508152 464636 508292 464656
rect 508112 464624 508158 464636
rect 502864 464532 502988 464542
rect 502864 464480 502874 464532
rect 502978 464526 502988 464532
rect 503088 464526 505668 464532
rect 505714 464530 505750 464620
rect 506092 464532 506216 464542
rect 502978 464492 503100 464526
rect 505656 464492 505668 464526
rect 502978 464480 502988 464492
rect 503088 464486 505668 464492
rect 502864 464470 502988 464480
rect 506092 464480 506102 464532
rect 506206 464516 506216 464532
rect 506280 464516 508080 464522
rect 506206 464482 506292 464516
rect 508068 464482 508080 464516
rect 506206 464480 506216 464482
rect 506092 464470 506216 464480
rect 506280 464476 508080 464482
rect 503088 464412 505668 464418
rect 503088 464378 503100 464412
rect 505656 464404 505668 464412
rect 505796 464412 506062 464418
rect 505796 464404 505802 464412
rect 505656 464378 505802 464404
rect 503088 464372 505802 464378
rect 505656 464370 505802 464372
rect 505796 464360 505802 464370
rect 506056 464404 506062 464412
rect 506280 464404 508080 464408
rect 506056 464402 508080 464404
rect 506056 464370 506292 464402
rect 506056 464360 506062 464370
rect 506280 464368 506292 464370
rect 508068 464368 508080 464402
rect 506280 464362 508080 464368
rect 505796 464354 506062 464360
rect 502606 464178 502738 464278
rect 505709 464268 505755 464270
rect 505702 464262 505772 464268
rect 505702 464054 505708 464262
rect 505766 464054 505772 464262
rect 505702 464048 505772 464054
rect 508112 464248 508158 464260
rect 508112 464064 508118 464248
rect 508152 464228 508432 464248
rect 508152 464084 508358 464228
rect 508412 464084 508432 464228
rect 508152 464064 508432 464084
rect 508112 464052 508158 464064
rect 502864 463960 502988 463970
rect 506092 463960 506216 463970
rect 502864 463908 502874 463960
rect 502978 463954 502988 463960
rect 503088 463954 505668 463960
rect 502978 463920 503100 463954
rect 505656 463920 505668 463954
rect 502978 463908 502988 463920
rect 503088 463914 505668 463920
rect 502864 463902 502988 463908
rect 506092 463908 506102 463960
rect 506206 463944 506216 463960
rect 506280 463944 508080 463950
rect 506206 463910 506292 463944
rect 508068 463910 508080 463944
rect 506206 463908 506216 463910
rect 506092 463898 506216 463908
rect 506280 463904 508080 463910
rect 500364 463810 501424 463850
rect 500364 463710 500398 463810
rect 500498 463710 500622 463810
rect 500722 463710 500846 463810
rect 500946 463710 501070 463810
rect 501170 463710 501294 463810
rect 501394 463710 501424 463810
rect 502664 463848 502788 463858
rect 502664 463796 502674 463848
rect 502778 463844 502788 463848
rect 503088 463844 505668 463846
rect 502778 463840 505668 463844
rect 502778 463806 503100 463840
rect 505656 463806 505668 463840
rect 502778 463802 505668 463806
rect 502778 463796 502788 463802
rect 503088 463800 505668 463802
rect 506280 463830 508158 463836
rect 502664 463786 502788 463796
rect 506280 463796 506292 463830
rect 508068 463796 508158 463830
rect 506280 463790 508158 463796
rect 500364 463586 501424 463710
rect 500364 463486 500398 463586
rect 500498 463486 500622 463586
rect 500722 463486 500846 463586
rect 500946 463486 501070 463586
rect 501170 463486 501294 463586
rect 501394 463486 501424 463586
rect 505708 463686 506062 463698
rect 505708 463502 505715 463686
rect 505749 463612 506062 463686
rect 505749 463560 505802 463612
rect 506056 463560 506062 463612
rect 505749 463502 506062 463560
rect 505708 463490 506062 463502
rect 508112 463676 508158 463790
rect 508112 463492 508118 463676
rect 508152 463492 508158 463676
rect 500364 463362 501424 463486
rect 500364 463262 500398 463362
rect 500498 463262 500622 463362
rect 500722 463262 500846 463362
rect 500946 463262 501070 463362
rect 501170 463262 501294 463362
rect 501394 463262 501424 463362
rect 502864 463388 502988 463398
rect 502864 463336 502874 463388
rect 502978 463382 502988 463388
rect 503088 463382 505668 463388
rect 502978 463348 503100 463382
rect 505656 463348 505668 463382
rect 508112 463378 508158 463492
rect 502978 463336 502988 463348
rect 503088 463342 505668 463348
rect 506280 463372 508158 463378
rect 502864 463330 502988 463336
rect 506280 463338 506292 463372
rect 508068 463338 508158 463372
rect 506280 463332 508158 463338
rect 500364 463138 501424 463262
rect 502664 463276 502788 463286
rect 502664 463224 502674 463276
rect 502778 463272 502788 463276
rect 503088 463272 505668 463274
rect 502778 463268 505668 463272
rect 502778 463234 503100 463268
rect 505656 463234 505668 463268
rect 502778 463230 505668 463234
rect 502778 463224 502788 463230
rect 503088 463228 505668 463230
rect 502664 463214 502788 463224
rect 500364 463038 500398 463138
rect 500498 463038 500622 463138
rect 500722 463038 500846 463138
rect 500946 463038 501070 463138
rect 501170 463038 501294 463138
rect 501394 463038 501424 463138
rect 500364 462914 501424 463038
rect 505708 463114 506062 463138
rect 505708 462930 505715 463114
rect 505749 463052 506062 463114
rect 505749 463000 505802 463052
rect 506056 463000 506062 463052
rect 505749 462930 506062 463000
rect 505709 462918 505755 462930
rect 500364 462814 500398 462914
rect 500498 462814 500622 462914
rect 500722 462814 500846 462914
rect 500946 462814 501070 462914
rect 501170 462814 501294 462914
rect 501394 462814 501424 462914
rect 506452 462894 508084 462902
rect 508112 462894 508158 463332
rect 506452 462886 508158 462894
rect 500364 462690 501424 462814
rect 502864 462816 502988 462826
rect 502864 462764 502874 462816
rect 502978 462810 502988 462816
rect 503088 462810 505668 462816
rect 502978 462776 503100 462810
rect 505656 462776 505668 462810
rect 502978 462764 502988 462776
rect 503088 462770 505668 462776
rect 506452 462786 506470 462886
rect 508068 462786 508158 462886
rect 506452 462780 508158 462786
rect 506452 462770 508084 462780
rect 502864 462758 502988 462764
rect 509464 462740 509786 468116
rect 509820 462740 509826 468116
rect 509464 462728 509826 462740
rect 510238 468116 510470 468128
rect 510238 462740 510244 468116
rect 510278 462740 510470 468116
rect 510238 462728 510470 462740
rect 500364 462590 500398 462690
rect 500498 462590 500622 462690
rect 500722 462590 500846 462690
rect 500946 462590 501070 462690
rect 501170 462590 501294 462690
rect 501394 462590 501424 462690
rect 502664 462704 502788 462714
rect 502664 462652 502674 462704
rect 502778 462700 502788 462704
rect 503088 462700 505668 462702
rect 502778 462696 505668 462700
rect 502778 462662 503100 462696
rect 505656 462662 505668 462696
rect 502778 462658 505668 462662
rect 502778 462652 502788 462658
rect 503088 462656 505668 462658
rect 502664 462642 502788 462652
rect 500364 462466 501424 462590
rect 509464 462578 509820 462728
rect 500364 462366 500398 462466
rect 500498 462366 500622 462466
rect 500722 462366 500846 462466
rect 500946 462366 501070 462466
rect 501170 462366 501294 462466
rect 501394 462366 501424 462466
rect 505708 462542 509820 462578
rect 505708 462370 505715 462542
rect 500364 462242 501424 462366
rect 505709 462358 505715 462370
rect 505749 462492 509820 462542
rect 505749 462440 505802 462492
rect 506056 462440 509820 462492
rect 505749 462370 509820 462440
rect 510258 462376 510470 462728
rect 510814 462376 510826 468840
rect 505749 462358 505755 462370
rect 510258 462364 510826 462376
rect 505709 462346 505755 462358
rect 500364 462142 500398 462242
rect 500498 462142 500622 462242
rect 500722 462142 500846 462242
rect 500946 462142 501070 462242
rect 501170 462142 501294 462242
rect 501394 462142 501424 462242
rect 502864 462244 502988 462254
rect 502864 462192 502874 462244
rect 502978 462238 502988 462244
rect 503088 462238 505668 462244
rect 502978 462204 503100 462238
rect 505656 462204 505668 462238
rect 502978 462192 502988 462204
rect 503088 462198 505668 462204
rect 502864 462186 502988 462192
rect 500364 462018 501424 462142
rect 502864 462134 502988 462144
rect 502864 462082 502874 462134
rect 502978 462130 502988 462134
rect 502978 462124 505756 462130
rect 502978 462090 503100 462124
rect 505656 462090 505756 462124
rect 502978 462084 505756 462090
rect 502978 462082 502988 462084
rect 502864 462072 502988 462082
rect 500364 461918 500398 462018
rect 500498 461918 500622 462018
rect 500722 461918 500846 462018
rect 500946 461918 501070 462018
rect 501170 461918 501294 462018
rect 501394 461918 501424 462018
rect 500364 461794 501424 461918
rect 500364 461694 500398 461794
rect 500498 461694 500622 461794
rect 500722 461694 500846 461794
rect 500946 461694 501070 461794
rect 501170 461694 501294 461794
rect 501394 461694 501424 461794
rect 500364 461570 501424 461694
rect 505708 461970 505756 462084
rect 505708 461786 505715 461970
rect 505749 461786 505756 461970
rect 502864 461676 502988 461686
rect 502864 461624 502874 461676
rect 502978 461672 502988 461676
rect 505708 461672 505756 461786
rect 502978 461666 505756 461672
rect 502978 461632 503100 461666
rect 505656 461632 505756 461666
rect 502978 461626 505756 461632
rect 502978 461624 502988 461626
rect 502864 461614 502988 461624
rect 500364 461470 500398 461570
rect 500498 461470 500622 461570
rect 500722 461470 500846 461570
rect 500946 461470 501070 461570
rect 501170 461470 501294 461570
rect 501394 461470 501424 461570
rect 500364 461346 501424 461470
rect 500364 461246 500398 461346
rect 500498 461246 500622 461346
rect 500722 461246 500846 461346
rect 500946 461246 501070 461346
rect 501170 461246 501294 461346
rect 501394 461246 501424 461346
rect 500364 461122 501424 461246
rect 508206 461310 512110 461316
rect 508206 461200 508212 461310
rect 508292 461200 511532 461310
rect 508206 461190 511532 461200
rect 511824 461190 512110 461310
rect 525660 461254 525666 472498
rect 526492 461254 526498 472498
rect 527584 472488 528644 472612
rect 527584 472388 527618 472488
rect 527718 472388 527842 472488
rect 527942 472388 528066 472488
rect 528166 472388 528290 472488
rect 528390 472388 528514 472488
rect 528614 472388 528644 472488
rect 527584 472264 528644 472388
rect 527584 472164 527618 472264
rect 527718 472164 527842 472264
rect 527942 472164 528066 472264
rect 528166 472164 528290 472264
rect 528390 472164 528514 472264
rect 528614 472164 528644 472264
rect 527584 472040 528644 472164
rect 527584 471940 527618 472040
rect 527718 471940 527842 472040
rect 527942 471940 528066 472040
rect 528166 471940 528290 472040
rect 528390 471940 528514 472040
rect 528614 471940 528644 472040
rect 527584 471816 528644 471940
rect 527584 471716 527618 471816
rect 527718 471716 527842 471816
rect 527942 471716 528066 471816
rect 528166 471716 528290 471816
rect 528390 471716 528514 471816
rect 528614 471716 528644 471816
rect 527584 471592 528644 471716
rect 527584 471492 527618 471592
rect 527718 471492 527842 471592
rect 527942 471492 528066 471592
rect 528166 471492 528290 471592
rect 528390 471492 528514 471592
rect 528614 471492 528644 471592
rect 527584 471368 528644 471492
rect 527584 471268 527618 471368
rect 527718 471268 527842 471368
rect 527942 471268 528066 471368
rect 528166 471268 528290 471368
rect 528390 471268 528514 471368
rect 528614 471268 528644 471368
rect 527584 471144 528644 471268
rect 527584 471044 527618 471144
rect 527718 471044 527842 471144
rect 527942 471044 528066 471144
rect 528166 471044 528290 471144
rect 528390 471044 528514 471144
rect 528614 471044 528644 471144
rect 527584 470920 528644 471044
rect 527584 470820 527618 470920
rect 527718 470820 527842 470920
rect 527942 470820 528066 470920
rect 528166 470820 528290 470920
rect 528390 470820 528514 470920
rect 528614 470820 528644 470920
rect 527584 470696 528644 470820
rect 527584 470596 527618 470696
rect 527718 470596 527842 470696
rect 527942 470596 528066 470696
rect 528166 470596 528290 470696
rect 528390 470596 528514 470696
rect 528614 470596 528644 470696
rect 527584 470472 528644 470596
rect 527584 470372 527618 470472
rect 527718 470372 527842 470472
rect 527942 470372 528066 470472
rect 528166 470372 528290 470472
rect 528390 470372 528514 470472
rect 528614 470372 528644 470472
rect 527584 470248 528644 470372
rect 527584 470148 527618 470248
rect 527718 470148 527842 470248
rect 527942 470148 528066 470248
rect 528166 470148 528290 470248
rect 528390 470148 528514 470248
rect 528614 470148 528644 470248
rect 527584 470024 528644 470148
rect 527584 469924 527618 470024
rect 527718 469924 527842 470024
rect 527942 469924 528066 470024
rect 528166 469924 528290 470024
rect 528390 469924 528514 470024
rect 528614 469924 528644 470024
rect 527584 469800 528644 469924
rect 527584 469700 527618 469800
rect 527718 469700 527842 469800
rect 527942 469700 528066 469800
rect 528166 469700 528290 469800
rect 528390 469700 528514 469800
rect 528614 469700 528644 469800
rect 527584 469576 528644 469700
rect 527584 469476 527618 469576
rect 527718 469476 527842 469576
rect 527942 469476 528066 469576
rect 528166 469476 528290 469576
rect 528390 469476 528514 469576
rect 528614 469476 528644 469576
rect 527584 469352 528644 469476
rect 527584 469252 527618 469352
rect 527718 469252 527842 469352
rect 527942 469252 528066 469352
rect 528166 469252 528290 469352
rect 528390 469252 528514 469352
rect 528614 469252 528644 469352
rect 527584 469128 528644 469252
rect 527584 469028 527618 469128
rect 527718 469028 527842 469128
rect 527942 469028 528066 469128
rect 528166 469028 528290 469128
rect 528390 469028 528514 469128
rect 528614 469028 528644 469128
rect 527584 468904 528644 469028
rect 527584 468804 527618 468904
rect 527718 468804 527842 468904
rect 527942 468804 528066 468904
rect 528166 468804 528290 468904
rect 528390 468804 528514 468904
rect 528614 468804 528644 468904
rect 527584 468680 528644 468804
rect 527584 468580 527618 468680
rect 527718 468580 527842 468680
rect 527942 468580 528066 468680
rect 528166 468580 528290 468680
rect 528390 468580 528514 468680
rect 528614 468580 528644 468680
rect 527584 468456 528644 468580
rect 527584 468356 527618 468456
rect 527718 468356 527842 468456
rect 527942 468356 528066 468456
rect 528166 468356 528290 468456
rect 528390 468356 528514 468456
rect 528614 468356 528644 468456
rect 527584 468232 528644 468356
rect 527584 468132 527618 468232
rect 527718 468132 527842 468232
rect 527942 468132 528066 468232
rect 528166 468132 528290 468232
rect 528390 468132 528514 468232
rect 528614 468132 528644 468232
rect 527584 468008 528644 468132
rect 527584 467908 527618 468008
rect 527718 467908 527842 468008
rect 527942 467908 528066 468008
rect 528166 467908 528290 468008
rect 528390 467908 528514 468008
rect 528614 467908 528644 468008
rect 527584 467784 528644 467908
rect 527584 467684 527618 467784
rect 527718 467684 527842 467784
rect 527942 467684 528066 467784
rect 528166 467684 528290 467784
rect 528390 467684 528514 467784
rect 528614 467684 528644 467784
rect 527584 467660 528644 467684
rect 525660 461248 526498 461254
rect 527584 463810 528644 463850
rect 527584 463710 527618 463810
rect 527718 463710 527842 463810
rect 527942 463710 528066 463810
rect 528166 463710 528290 463810
rect 528390 463710 528514 463810
rect 528614 463710 528644 463810
rect 527584 463586 528644 463710
rect 527584 463486 527618 463586
rect 527718 463486 527842 463586
rect 527942 463486 528066 463586
rect 528166 463486 528290 463586
rect 528390 463486 528514 463586
rect 528614 463486 528644 463586
rect 527584 463362 528644 463486
rect 527584 463262 527618 463362
rect 527718 463262 527842 463362
rect 527942 463262 528066 463362
rect 528166 463262 528290 463362
rect 528390 463262 528514 463362
rect 528614 463262 528644 463362
rect 527584 463138 528644 463262
rect 527584 463038 527618 463138
rect 527718 463038 527842 463138
rect 527942 463038 528066 463138
rect 528166 463038 528290 463138
rect 528390 463038 528514 463138
rect 528614 463038 528644 463138
rect 527584 462914 528644 463038
rect 527584 462814 527618 462914
rect 527718 462814 527842 462914
rect 527942 462814 528066 462914
rect 528166 462814 528290 462914
rect 528390 462814 528514 462914
rect 528614 462814 528644 462914
rect 527584 462690 528644 462814
rect 527584 462590 527618 462690
rect 527718 462590 527842 462690
rect 527942 462590 528066 462690
rect 528166 462590 528290 462690
rect 528390 462590 528514 462690
rect 528614 462590 528644 462690
rect 527584 462466 528644 462590
rect 527584 462366 527618 462466
rect 527718 462366 527842 462466
rect 527942 462366 528066 462466
rect 528166 462366 528290 462466
rect 528390 462366 528514 462466
rect 528614 462366 528644 462466
rect 527584 462242 528644 462366
rect 527584 462142 527618 462242
rect 527718 462142 527842 462242
rect 527942 462142 528066 462242
rect 528166 462142 528290 462242
rect 528390 462142 528514 462242
rect 528614 462142 528644 462242
rect 527584 462018 528644 462142
rect 527584 461918 527618 462018
rect 527718 461918 527842 462018
rect 527942 461918 528066 462018
rect 528166 461918 528290 462018
rect 528390 461918 528514 462018
rect 528614 461918 528644 462018
rect 527584 461794 528644 461918
rect 527584 461694 527618 461794
rect 527718 461694 527842 461794
rect 527942 461694 528066 461794
rect 528166 461694 528290 461794
rect 528390 461694 528514 461794
rect 528614 461694 528644 461794
rect 527584 461570 528644 461694
rect 527584 461470 527618 461570
rect 527718 461470 527842 461570
rect 527942 461470 528066 461570
rect 528166 461470 528290 461570
rect 528390 461470 528514 461570
rect 528614 461470 528644 461570
rect 527584 461346 528644 461470
rect 508206 461184 512110 461190
rect 527584 461246 527618 461346
rect 527718 461246 527842 461346
rect 527942 461246 528066 461346
rect 528166 461246 528290 461346
rect 528390 461246 528514 461346
rect 528614 461246 528644 461346
rect 500364 461022 500398 461122
rect 500498 461022 500622 461122
rect 500722 461022 500846 461122
rect 500946 461022 501070 461122
rect 501170 461022 501294 461122
rect 501394 461022 501424 461122
rect 527584 461122 528644 461246
rect 500364 460898 501424 461022
rect 502864 461074 505580 461090
rect 502864 461064 503226 461074
rect 502864 461012 502874 461064
rect 502978 461012 503226 461064
rect 502864 460974 503226 461012
rect 505568 460974 505580 461074
rect 502864 460958 505580 460974
rect 527584 461022 527618 461122
rect 527718 461022 527842 461122
rect 527942 461022 528066 461122
rect 528166 461022 528290 461122
rect 528390 461022 528514 461122
rect 528614 461022 528644 461122
rect 500364 460798 500398 460898
rect 500498 460798 500622 460898
rect 500722 460798 500846 460898
rect 500946 460798 501070 460898
rect 501170 460798 501294 460898
rect 501394 460798 501424 460898
rect 527584 460898 528644 461022
rect 500364 460674 501424 460798
rect 508346 460854 512536 460860
rect 508346 460734 508352 460854
rect 508432 460734 512116 460854
rect 512530 460734 512536 460854
rect 508346 460728 512536 460734
rect 527584 460798 527618 460898
rect 527718 460798 527842 460898
rect 527942 460798 528066 460898
rect 528166 460798 528290 460898
rect 528390 460798 528514 460898
rect 528614 460798 528644 460898
rect 500364 460574 500398 460674
rect 500498 460574 500622 460674
rect 500722 460574 500846 460674
rect 500946 460574 501070 460674
rect 501170 460574 501294 460674
rect 501394 460574 501424 460674
rect 500364 460450 501424 460574
rect 527584 460674 528644 460798
rect 527584 460574 527618 460674
rect 527718 460574 527842 460674
rect 527942 460574 528066 460674
rect 528166 460574 528290 460674
rect 528390 460574 528514 460674
rect 528614 460574 528644 460674
rect 500364 460350 500398 460450
rect 500498 460350 500622 460450
rect 500722 460350 500846 460450
rect 500946 460350 501070 460450
rect 501170 460350 501294 460450
rect 501394 460350 501424 460450
rect 500364 460226 501424 460350
rect 500364 460126 500398 460226
rect 500498 460126 500622 460226
rect 500722 460126 500846 460226
rect 500946 460126 501070 460226
rect 501170 460126 501294 460226
rect 501394 460126 501424 460226
rect 500364 460002 501424 460126
rect 500364 459902 500398 460002
rect 500498 459902 500622 460002
rect 500722 459902 500846 460002
rect 500946 459902 501070 460002
rect 501170 459902 501294 460002
rect 501394 459902 501424 460002
rect 500364 459778 501424 459902
rect 500364 459678 500398 459778
rect 500498 459678 500622 459778
rect 500722 459678 500846 459778
rect 500946 459678 501070 459778
rect 501170 459678 501294 459778
rect 501394 459678 501424 459778
rect 500364 459554 501424 459678
rect 500364 459454 500398 459554
rect 500498 459454 500622 459554
rect 500722 459454 500846 459554
rect 500946 459454 501070 459554
rect 501170 459454 501294 459554
rect 501394 459454 501424 459554
rect 500364 459330 501424 459454
rect 500364 459230 500398 459330
rect 500498 459230 500622 459330
rect 500722 459230 500846 459330
rect 500946 459230 501070 459330
rect 501170 459230 501294 459330
rect 501394 459230 501424 459330
rect 502428 460352 502728 460452
rect 527584 460450 528644 460574
rect 502428 459952 502528 460352
rect 502628 459952 502728 460352
rect 502808 460442 506062 460448
rect 502808 459974 502814 460442
rect 502962 459974 505802 460442
rect 506056 459974 506062 460442
rect 502808 459968 506062 459974
rect 527584 460350 527618 460450
rect 527718 460350 527842 460450
rect 527942 460350 528066 460450
rect 528166 460350 528290 460450
rect 528390 460350 528514 460450
rect 528614 460350 528644 460450
rect 527584 460226 528644 460350
rect 527584 460126 527618 460226
rect 527718 460126 527842 460226
rect 527942 460126 528066 460226
rect 528166 460126 528290 460226
rect 528390 460126 528514 460226
rect 528614 460126 528644 460226
rect 527584 460002 528644 460126
rect 502428 459758 502728 459952
rect 527584 459902 527618 460002
rect 527718 459902 527842 460002
rect 527942 459902 528066 460002
rect 528166 459902 528290 460002
rect 528390 459902 528514 460002
rect 528614 459902 528644 460002
rect 517858 459868 518267 459880
rect 502428 459752 510866 459758
rect 502428 459718 503138 459752
rect 510854 459718 510866 459752
rect 502428 459712 510866 459718
rect 502428 459610 503086 459712
rect 502428 459598 503085 459610
rect 502428 459414 503045 459598
rect 503079 459418 503085 459598
rect 503079 459414 503086 459418
rect 502428 459300 503086 459414
rect 510928 459336 513328 459342
rect 510928 459302 512134 459336
rect 510828 459300 512134 459302
rect 503122 459294 512134 459300
rect 503122 459260 503138 459294
rect 510854 459262 512134 459294
rect 510854 459260 510866 459262
rect 503122 459254 510866 459260
rect 500364 459106 501424 459230
rect 503039 459142 503085 459152
rect 500364 459006 500398 459106
rect 500498 459006 500622 459106
rect 500722 459006 500846 459106
rect 500946 459006 501070 459106
rect 501170 459006 501294 459106
rect 501394 459006 501424 459106
rect 500364 458882 501424 459006
rect 502808 459140 503088 459142
rect 502808 459122 503045 459140
rect 502808 458982 502828 459122
rect 502948 458982 503045 459122
rect 502808 458962 503045 458982
rect 503039 458956 503045 458962
rect 503079 458962 503088 459140
rect 503079 458956 503085 458962
rect 503039 458944 503085 458956
rect 500364 458782 500398 458882
rect 500498 458782 500622 458882
rect 500722 458782 500846 458882
rect 500946 458782 501070 458882
rect 501170 458782 501294 458882
rect 501394 458782 501424 458882
rect 500364 458658 501424 458782
rect 502648 458862 502768 458882
rect 502648 458782 502668 458862
rect 502748 458842 502768 458862
rect 502748 458836 510866 458842
rect 502748 458802 503138 458836
rect 510854 458802 510866 458836
rect 502748 458782 502768 458802
rect 503126 458796 510866 458802
rect 502648 458762 502768 458782
rect 503039 458682 503085 458694
rect 500364 458558 500398 458658
rect 500498 458558 500622 458658
rect 500722 458558 500846 458658
rect 500946 458558 501070 458658
rect 501170 458558 501294 458658
rect 501394 458558 501424 458658
rect 500364 458434 501424 458558
rect 502808 458662 503045 458682
rect 502808 458522 502828 458662
rect 502948 458522 503045 458662
rect 502808 458502 503045 458522
rect 503039 458498 503045 458502
rect 503079 458502 503088 458682
rect 503079 458498 503085 458502
rect 503039 458486 503085 458498
rect 500364 458334 500398 458434
rect 500498 458334 500622 458434
rect 500722 458334 500846 458434
rect 500946 458334 501070 458434
rect 501170 458334 501294 458434
rect 501394 458334 501424 458434
rect 503126 458382 510866 458384
rect 510928 458382 512134 459262
rect 503126 458378 512134 458382
rect 503126 458344 503138 458378
rect 510854 458344 512134 458378
rect 503126 458342 512134 458344
rect 503126 458338 510866 458342
rect 500364 458210 501424 458334
rect 503039 458224 503085 458236
rect 503039 458222 503045 458224
rect 500364 458110 500398 458210
rect 500498 458110 500622 458210
rect 500722 458110 500846 458210
rect 500946 458110 501070 458210
rect 501170 458110 501294 458210
rect 501394 458110 501424 458210
rect 500364 457986 501424 458110
rect 502808 458202 503045 458222
rect 502808 458062 502828 458202
rect 502948 458062 503045 458202
rect 502808 458042 503045 458062
rect 503039 458040 503045 458042
rect 503079 458222 503085 458224
rect 503079 458042 503088 458222
rect 503079 458040 503085 458042
rect 503039 458028 503085 458040
rect 500364 457886 500398 457986
rect 500498 457886 500622 457986
rect 500722 457886 500846 457986
rect 500946 457886 501070 457986
rect 501170 457886 501294 457986
rect 501394 457886 501424 457986
rect 500364 457762 501424 457886
rect 502648 457942 502768 457962
rect 502648 457862 502668 457942
rect 502748 457922 502768 457942
rect 503126 457922 510866 457926
rect 502748 457920 510866 457922
rect 502748 457886 503138 457920
rect 510854 457886 510866 457920
rect 502748 457882 510866 457886
rect 502748 457862 502768 457882
rect 503126 457880 510866 457882
rect 502648 457842 502768 457862
rect 503039 457766 503085 457778
rect 503039 457762 503045 457766
rect 500364 457662 500398 457762
rect 500498 457662 500622 457762
rect 500722 457662 500846 457762
rect 500946 457662 501070 457762
rect 501170 457662 501294 457762
rect 501394 457662 501424 457762
rect 500364 457538 501424 457662
rect 502808 457742 503045 457762
rect 502808 457602 502828 457742
rect 502948 457602 503045 457742
rect 502808 457582 503045 457602
rect 503079 457762 503085 457766
rect 503079 457582 503088 457762
rect 503039 457570 503085 457582
rect 500364 457438 500398 457538
rect 500498 457438 500622 457538
rect 500722 457438 500846 457538
rect 500946 457438 501070 457538
rect 501170 457438 501294 457538
rect 501394 457438 501424 457538
rect 500364 457314 501424 457438
rect 503126 457462 510866 457468
rect 510928 457462 512134 458342
rect 503126 457428 503138 457462
rect 510854 457428 512134 457462
rect 503126 457422 512134 457428
rect 510928 457348 512134 457422
rect 512422 457348 512836 459336
rect 513286 457348 513328 459336
rect 517858 459330 517864 459868
rect 518261 459330 518267 459868
rect 517858 459318 518267 459330
rect 521613 459868 522022 459880
rect 521613 459330 521619 459868
rect 522016 459330 522022 459868
rect 521613 459318 522022 459330
rect 527584 459778 528644 459902
rect 527584 459678 527618 459778
rect 527718 459678 527842 459778
rect 527942 459678 528066 459778
rect 528166 459678 528290 459778
rect 528390 459678 528514 459778
rect 528614 459678 528644 459778
rect 527584 459554 528644 459678
rect 527584 459454 527618 459554
rect 527718 459454 527842 459554
rect 527942 459454 528066 459554
rect 528166 459454 528290 459554
rect 528390 459454 528514 459554
rect 528614 459454 528644 459554
rect 527584 459330 528644 459454
rect 527584 459230 527618 459330
rect 527718 459230 527842 459330
rect 527942 459230 528066 459330
rect 528166 459230 528290 459330
rect 528390 459230 528514 459330
rect 528614 459230 528644 459330
rect 527584 459106 528644 459230
rect 510928 457342 513328 457348
rect 516852 459050 518278 459066
rect 516852 458512 517864 459050
rect 518261 458512 518278 459050
rect 516852 458496 518278 458512
rect 521613 459050 522022 459062
rect 521613 458512 521619 459050
rect 522016 458512 522022 459050
rect 521613 458500 522022 458512
rect 527584 459006 527618 459106
rect 527718 459006 527842 459106
rect 527942 459006 528066 459106
rect 528166 459006 528290 459106
rect 528390 459006 528514 459106
rect 528614 459006 528644 459106
rect 527584 458882 528644 459006
rect 527584 458782 527618 458882
rect 527718 458782 527842 458882
rect 527942 458782 528066 458882
rect 528166 458782 528290 458882
rect 528390 458782 528514 458882
rect 528614 458782 528644 458882
rect 527584 458658 528644 458782
rect 527584 458558 527618 458658
rect 527718 458558 527842 458658
rect 527942 458558 528066 458658
rect 528166 458558 528290 458658
rect 528390 458558 528514 458658
rect 528614 458558 528644 458658
rect 500364 457214 500398 457314
rect 500498 457214 500622 457314
rect 500722 457214 500846 457314
rect 500946 457214 501070 457314
rect 501170 457214 501294 457314
rect 501394 457214 501424 457314
rect 503039 457308 503085 457320
rect 503039 457302 503045 457308
rect 500364 457190 501424 457214
rect 502808 457282 503045 457302
rect 502808 457142 502828 457282
rect 502948 457142 503045 457282
rect 502808 457124 503045 457142
rect 503079 457302 503085 457308
rect 503079 457124 503088 457302
rect 502808 457122 503088 457124
rect 503039 457112 503085 457122
rect 502648 457022 502768 457042
rect 502648 456942 502668 457022
rect 502748 457002 502768 457022
rect 503126 457004 510866 457010
rect 503126 457002 503138 457004
rect 502748 456970 503138 457002
rect 510854 456970 510866 457004
rect 502748 456964 510866 456970
rect 502748 456962 503148 456964
rect 502748 456942 502768 456962
rect 502648 456922 502768 456942
rect 503039 456850 503085 456862
rect 503039 456842 503045 456850
rect 502808 456822 503045 456842
rect 502808 456682 502828 456822
rect 502948 456682 503045 456822
rect 502808 456666 503045 456682
rect 503079 456842 503085 456850
rect 503079 456666 503088 456842
rect 502808 456662 503088 456666
rect 503039 456654 503085 456662
rect 510928 456636 511834 456642
rect 510928 456562 511534 456636
rect 510848 456552 511534 456562
rect 503126 456546 511534 456552
rect 503126 456512 503138 456546
rect 510854 456512 511534 456546
rect 503126 456506 511534 456512
rect 510848 456502 511534 456506
rect 503039 456392 503085 456404
rect 503039 456382 503045 456392
rect 502808 456362 503045 456382
rect 502808 456222 502828 456362
rect 502948 456222 503045 456362
rect 502808 456208 503045 456222
rect 503079 456382 503085 456392
rect 503079 456208 503088 456382
rect 502808 456202 503088 456208
rect 503039 456196 503085 456202
rect 502648 456102 502768 456122
rect 502648 456022 502668 456102
rect 502748 456094 503148 456102
rect 502748 456088 510866 456094
rect 502748 456062 503138 456088
rect 502748 456022 502768 456062
rect 503126 456054 503138 456062
rect 510854 456054 510866 456088
rect 503126 456048 510866 456054
rect 502648 456002 502768 456022
rect 503039 455934 503085 455946
rect 503039 455922 503045 455934
rect 502808 455902 503045 455922
rect 502808 455762 502828 455902
rect 502948 455762 503045 455902
rect 502808 455750 503045 455762
rect 503079 455922 503085 455934
rect 503079 455750 503088 455922
rect 502808 455742 503088 455750
rect 503039 455738 503085 455742
rect 510928 455642 511534 456502
rect 510828 455636 511534 455642
rect 503126 455630 511534 455636
rect 503126 455596 503138 455630
rect 510854 455596 511534 455630
rect 503126 455590 511534 455596
rect 510828 455582 511534 455590
rect 503039 455476 503085 455488
rect 503039 455462 503045 455476
rect 502808 455442 503045 455462
rect 502808 455302 502828 455442
rect 502948 455302 503045 455442
rect 502808 455292 503045 455302
rect 503079 455462 503085 455476
rect 503079 455292 503088 455462
rect 502808 455282 503088 455292
rect 503039 455280 503085 455282
rect 502648 455182 502768 455202
rect 502648 455102 502668 455182
rect 502748 455178 503148 455182
rect 502748 455172 510866 455178
rect 502748 455142 503138 455172
rect 502748 455102 502768 455142
rect 503126 455138 503138 455142
rect 510854 455138 510866 455172
rect 503126 455132 510866 455138
rect 502648 455082 502768 455102
rect 503039 455018 503085 455030
rect 503039 455002 503045 455018
rect 502808 454982 503045 455002
rect 502808 454842 502828 454982
rect 502948 454842 503045 454982
rect 502808 454834 503045 454842
rect 503079 455002 503085 455018
rect 503079 454834 503088 455002
rect 502808 454822 503088 454834
rect 510928 454722 511534 455582
rect 510828 454720 511534 454722
rect 503126 454714 511534 454720
rect 503126 454680 503138 454714
rect 510854 454680 511534 454714
rect 503126 454674 511534 454680
rect 510828 454662 511534 454674
rect 510928 454648 511534 454662
rect 511822 454648 511834 456636
rect 510928 454642 511834 454648
rect 502428 454442 502728 454542
rect 502428 454042 502528 454442
rect 502628 454042 502728 454442
rect 502428 453942 502728 454042
rect 510926 453802 514926 453842
rect 510848 453800 514926 453802
rect 503126 453794 514926 453800
rect 503126 453760 503138 453794
rect 510854 453762 514926 453794
rect 510854 453760 510866 453762
rect 503126 453754 510866 453760
rect 510926 453756 514926 453762
rect 503039 453642 503085 453652
rect 502808 453640 503088 453642
rect 502808 453622 503045 453640
rect 502808 453482 502828 453622
rect 502948 453482 503045 453622
rect 502808 453462 503045 453482
rect 503039 453456 503045 453462
rect 503079 453462 503088 453640
rect 510926 453556 513720 453756
rect 513920 453556 514154 453756
rect 514354 453556 514588 453756
rect 514788 453556 514926 453756
rect 503079 453456 503085 453462
rect 503039 453444 503085 453456
rect 502648 453362 502768 453382
rect 502648 453282 502668 453362
rect 502748 453342 502768 453362
rect 502748 453336 510866 453342
rect 502748 453302 503138 453336
rect 510854 453302 510866 453336
rect 502748 453282 502768 453302
rect 503126 453296 510866 453302
rect 510926 453322 514926 453556
rect 502648 453262 502768 453282
rect 503039 453182 503085 453194
rect 502808 453162 503045 453182
rect 502808 453022 502828 453162
rect 502948 453022 503045 453162
rect 502808 453002 503045 453022
rect 503039 452998 503045 453002
rect 503079 453002 503088 453182
rect 510926 453122 513720 453322
rect 513920 453122 514154 453322
rect 514354 453122 514588 453322
rect 514788 453122 514926 453322
rect 503079 452998 503085 453002
rect 503039 452986 503085 452998
rect 510926 452888 514926 453122
rect 503126 452882 510866 452884
rect 510926 452882 513720 452888
rect 503126 452878 513720 452882
rect 503126 452844 503138 452878
rect 510854 452844 513720 452878
rect 503126 452842 513720 452844
rect 503126 452838 510866 452842
rect 503039 452724 503085 452736
rect 503039 452722 503045 452724
rect 502808 452702 503045 452722
rect 502808 452562 502828 452702
rect 502948 452562 503045 452702
rect 502808 452542 503045 452562
rect 503039 452540 503045 452542
rect 503079 452722 503085 452724
rect 503079 452542 503088 452722
rect 510926 452688 513720 452842
rect 513920 452688 514154 452888
rect 514354 452688 514588 452888
rect 514788 452688 514926 452888
rect 503079 452540 503085 452542
rect 503039 452528 503085 452540
rect 502648 452442 502768 452462
rect 502648 452362 502668 452442
rect 502748 452422 502768 452442
rect 510926 452454 514926 452688
rect 503126 452422 510866 452426
rect 502748 452420 510866 452422
rect 502748 452386 503138 452420
rect 510854 452386 510866 452420
rect 502748 452382 510866 452386
rect 502748 452362 502768 452382
rect 503126 452380 510866 452382
rect 502648 452342 502768 452362
rect 503039 452266 503085 452278
rect 503039 452262 503045 452266
rect 502808 452242 503045 452262
rect 502808 452102 502828 452242
rect 502948 452102 503045 452242
rect 502808 452082 503045 452102
rect 503079 452262 503085 452266
rect 503079 452082 503088 452262
rect 510926 452254 513720 452454
rect 513920 452254 514154 452454
rect 514354 452254 514588 452454
rect 514788 452254 514926 452454
rect 503039 452070 503085 452082
rect 510926 452020 514926 452254
rect 503126 451962 510866 451968
rect 510926 451962 513720 452020
rect 503126 451928 503138 451962
rect 510854 451928 513720 451962
rect 503126 451922 513720 451928
rect 510926 451820 513720 451922
rect 513920 451820 514154 452020
rect 514354 451820 514588 452020
rect 514788 451820 514926 452020
rect 503039 451808 503085 451820
rect 503039 451802 503045 451808
rect 502808 451782 503045 451802
rect 502808 451642 502828 451782
rect 502948 451642 503045 451782
rect 502808 451624 503045 451642
rect 503079 451802 503085 451808
rect 503079 451624 503088 451802
rect 502808 451622 503088 451624
rect 503039 451612 503085 451622
rect 510926 451586 514926 451820
rect 502648 451522 502768 451542
rect 502648 451442 502668 451522
rect 502748 451502 502768 451522
rect 503126 451504 510866 451510
rect 503126 451502 503138 451504
rect 502748 451470 503138 451502
rect 510854 451470 510866 451504
rect 502748 451464 510866 451470
rect 502748 451462 503148 451464
rect 502748 451442 502768 451462
rect 502648 451422 502768 451442
rect 510926 451386 513720 451586
rect 513920 451386 514154 451586
rect 514354 451386 514588 451586
rect 514788 451386 514926 451586
rect 503039 451350 503085 451362
rect 503039 451342 503045 451350
rect 502808 451322 503045 451342
rect 502808 451182 502828 451322
rect 502948 451182 503045 451322
rect 502808 451166 503045 451182
rect 503079 451342 503085 451350
rect 503079 451166 503088 451342
rect 502808 451162 503088 451166
rect 503039 451154 503085 451162
rect 510926 451152 514926 451386
rect 503126 451046 510866 451052
rect 503126 451012 503138 451046
rect 510854 451042 510866 451046
rect 510926 451042 513720 451152
rect 510854 451012 513720 451042
rect 503126 451006 513720 451012
rect 510828 451002 513720 451006
rect 510926 450952 513720 451002
rect 513920 450952 514154 451152
rect 514354 450952 514588 451152
rect 514788 450952 514926 451152
rect 516202 451688 516611 451700
rect 516202 451150 516208 451688
rect 516605 451150 516611 451688
rect 516202 451138 516611 451150
rect 503039 450892 503085 450904
rect 503039 450882 503045 450892
rect 502808 450862 503045 450882
rect 502808 450722 502828 450862
rect 502948 450722 503045 450862
rect 502808 450708 503045 450722
rect 503079 450882 503085 450892
rect 503079 450708 503088 450882
rect 502808 450702 503088 450708
rect 510926 450718 514926 450952
rect 503039 450696 503085 450702
rect 502648 450602 502768 450622
rect 502648 450522 502668 450602
rect 502748 450594 503148 450602
rect 502748 450588 510866 450594
rect 502748 450562 503138 450588
rect 502748 450522 502768 450562
rect 503126 450554 503138 450562
rect 510854 450554 510866 450588
rect 503126 450548 510866 450554
rect 502648 450502 502768 450522
rect 510926 450518 513720 450718
rect 513920 450518 514154 450718
rect 514354 450518 514588 450718
rect 514788 450518 514926 450718
rect 503039 450434 503085 450446
rect 503039 450422 503045 450434
rect 502808 450402 503045 450422
rect 502808 450262 502828 450402
rect 502948 450262 503045 450402
rect 502808 450250 503045 450262
rect 503079 450422 503085 450434
rect 503079 450250 503088 450422
rect 502808 450242 503088 450250
rect 510926 450284 514926 450518
rect 503039 450238 503085 450242
rect 510926 450142 513720 450284
rect 510828 450136 513720 450142
rect 503126 450130 513720 450136
rect 503126 450096 503138 450130
rect 510854 450096 513720 450130
rect 503126 450090 513720 450096
rect 510828 450084 513720 450090
rect 513920 450084 514154 450284
rect 514354 450084 514588 450284
rect 514788 450084 514926 450284
rect 510828 450082 514926 450084
rect 503039 449976 503085 449988
rect 503039 449962 503045 449976
rect 502808 449942 503045 449962
rect 502808 449802 502828 449942
rect 502948 449802 503045 449942
rect 502808 449792 503045 449802
rect 503079 449962 503085 449976
rect 503079 449792 503088 449962
rect 502808 449782 503088 449792
rect 510926 449850 514926 450082
rect 503039 449780 503085 449782
rect 502648 449682 502768 449702
rect 502648 449602 502668 449682
rect 502748 449678 503148 449682
rect 502748 449672 510866 449678
rect 502748 449642 503138 449672
rect 502748 449602 502768 449642
rect 503126 449638 503138 449642
rect 510854 449638 510866 449672
rect 503126 449632 510866 449638
rect 510926 449650 513720 449850
rect 513920 449650 514154 449850
rect 514354 449650 514588 449850
rect 514788 449650 514926 449850
rect 502648 449582 502768 449602
rect 503039 449518 503085 449530
rect 503039 449502 503045 449518
rect 502808 449482 503045 449502
rect 502808 449342 502828 449482
rect 502948 449342 503045 449482
rect 502808 449334 503045 449342
rect 503079 449502 503085 449518
rect 503079 449334 503088 449502
rect 502808 449322 503088 449334
rect 510926 449416 514926 449650
rect 510926 449222 513720 449416
rect 510828 449220 513720 449222
rect 503126 449216 513720 449220
rect 513920 449216 514154 449416
rect 514354 449216 514588 449416
rect 514788 449216 514926 449416
rect 503126 449214 514926 449216
rect 503126 449180 503138 449214
rect 510854 449180 514926 449214
rect 503126 449174 514926 449180
rect 510828 449162 514926 449174
rect 510926 449142 514926 449162
rect 502428 448942 502728 449042
rect 502428 448542 502528 448942
rect 502628 448542 502728 448942
rect 502428 448442 502728 448542
rect 514234 449016 514926 449142
rect 514234 448816 514588 449016
rect 514788 448816 514926 449016
rect 514234 448616 514926 448816
rect 514234 448416 514588 448616
rect 514788 448416 514926 448616
rect 510928 448336 511834 448342
rect 510928 448302 511534 448336
rect 510828 448300 511534 448302
rect 503126 448294 511534 448300
rect 503126 448260 503138 448294
rect 510854 448262 511534 448294
rect 510854 448260 510866 448262
rect 503126 448254 510866 448260
rect 503039 448142 503085 448152
rect 502808 448140 503088 448142
rect 502808 448122 503045 448140
rect 502808 447982 502828 448122
rect 502948 447982 503045 448122
rect 502808 447962 503045 447982
rect 503039 447956 503045 447962
rect 503079 447962 503088 448140
rect 503079 447956 503085 447962
rect 503039 447944 503085 447956
rect 502648 447862 502768 447882
rect 502648 447782 502668 447862
rect 502748 447842 502768 447862
rect 502748 447836 510866 447842
rect 502748 447802 503138 447836
rect 510854 447802 510866 447836
rect 502748 447782 502768 447802
rect 503126 447796 510866 447802
rect 502648 447762 502768 447782
rect 503039 447682 503085 447694
rect 502808 447662 503045 447682
rect 502808 447522 502828 447662
rect 502948 447522 503045 447662
rect 502808 447502 503045 447522
rect 503039 447498 503045 447502
rect 503079 447502 503088 447682
rect 503079 447498 503085 447502
rect 503039 447486 503085 447498
rect 503126 447382 510866 447384
rect 510928 447382 511534 448262
rect 503126 447378 511534 447382
rect 503126 447344 503138 447378
rect 510854 447344 511534 447378
rect 503126 447342 511534 447344
rect 503126 447338 510866 447342
rect 503039 447224 503085 447236
rect 503039 447222 503045 447224
rect 502808 447202 503045 447222
rect 502808 447062 502828 447202
rect 502948 447062 503045 447202
rect 502808 447042 503045 447062
rect 503039 447040 503045 447042
rect 503079 447222 503085 447224
rect 503079 447042 503088 447222
rect 503079 447040 503085 447042
rect 503039 447028 503085 447040
rect 502648 446942 502768 446962
rect 502648 446862 502668 446942
rect 502748 446922 502768 446942
rect 503126 446922 510866 446926
rect 502748 446920 510866 446922
rect 502748 446886 503138 446920
rect 510854 446886 510866 446920
rect 502748 446882 510866 446886
rect 502748 446862 502768 446882
rect 503126 446880 510866 446882
rect 502648 446842 502768 446862
rect 503039 446766 503085 446778
rect 503039 446762 503045 446766
rect 502808 446742 503045 446762
rect 502808 446602 502828 446742
rect 502948 446602 503045 446742
rect 502808 446582 503045 446602
rect 503079 446762 503085 446766
rect 503079 446582 503088 446762
rect 503039 446570 503085 446582
rect 503126 446462 510866 446468
rect 510928 446462 511534 447342
rect 503126 446428 503138 446462
rect 510854 446428 511534 446462
rect 503126 446422 511534 446428
rect 510928 446348 511534 446422
rect 511822 446348 511834 448336
rect 510928 446342 511834 446348
rect 514234 448216 514926 448416
rect 514234 448016 514588 448216
rect 514788 448016 514926 448216
rect 514234 447816 514926 448016
rect 515390 450880 515960 450886
rect 515390 450322 515396 450880
rect 515954 450322 515960 450880
rect 515390 448426 515960 450322
rect 516190 450880 516622 450886
rect 516190 450322 516196 450880
rect 516616 450322 516622 450880
rect 516190 450316 516622 450322
rect 516190 450062 516622 450068
rect 516190 449504 516196 450062
rect 516616 449504 516622 450062
rect 516190 449498 516622 449504
rect 516190 449244 516622 449250
rect 516190 448686 516196 449244
rect 516616 448686 516622 449244
rect 516190 448680 516622 448686
rect 516852 449244 517422 458496
rect 527584 458434 528644 458558
rect 527584 458334 527618 458434
rect 527718 458334 527842 458434
rect 527942 458334 528066 458434
rect 528166 458334 528290 458434
rect 528390 458334 528514 458434
rect 528614 458334 528644 458434
rect 517858 458232 518267 458244
rect 517858 457694 517864 458232
rect 518261 457694 518267 458232
rect 517858 457682 518267 457694
rect 521613 458232 522022 458244
rect 521613 457694 521619 458232
rect 522016 457694 522022 458232
rect 521613 457682 522022 457694
rect 527584 458210 528644 458334
rect 527584 458110 527618 458210
rect 527718 458110 527842 458210
rect 527942 458110 528066 458210
rect 528166 458110 528290 458210
rect 528390 458110 528514 458210
rect 528614 458110 528644 458210
rect 527584 457986 528644 458110
rect 527584 457886 527618 457986
rect 527718 457886 527842 457986
rect 527942 457886 528066 457986
rect 528166 457886 528290 457986
rect 528390 457886 528514 457986
rect 528614 457886 528644 457986
rect 527584 457762 528644 457886
rect 527584 457662 527618 457762
rect 527718 457662 527842 457762
rect 527942 457662 528066 457762
rect 528166 457662 528290 457762
rect 528390 457662 528514 457762
rect 528614 457662 528644 457762
rect 527584 457538 528644 457662
rect 527584 457438 527618 457538
rect 527718 457438 527842 457538
rect 527942 457438 528066 457538
rect 528166 457438 528290 457538
rect 528390 457438 528514 457538
rect 528614 457438 528644 457538
rect 517552 457412 518688 457434
rect 517552 456918 517594 457412
rect 518660 456918 518688 457412
rect 527584 457314 528644 457438
rect 527584 457214 527618 457314
rect 527718 457214 527842 457314
rect 527942 457214 528066 457314
rect 528166 457214 528290 457314
rect 528390 457214 528514 457314
rect 528614 457214 528644 457314
rect 527584 457190 528644 457214
rect 517552 456596 518688 456918
rect 517552 456058 518274 456596
rect 518671 456058 518688 456596
rect 517552 455778 518688 456058
rect 522999 456596 523408 456608
rect 522999 456058 523005 456596
rect 523402 456058 523408 456596
rect 522999 456046 523408 456058
rect 517552 455240 518274 455778
rect 518671 455240 518688 455778
rect 517552 454960 518688 455240
rect 522988 455788 523420 455794
rect 522988 455230 522994 455788
rect 523414 455230 523420 455788
rect 522988 455224 523420 455230
rect 523588 455788 524158 455794
rect 523588 455230 523594 455788
rect 524152 455230 524158 455788
rect 517552 454422 518274 454960
rect 518671 454422 518688 454960
rect 517552 454142 518688 454422
rect 517552 453604 518274 454142
rect 518671 453604 518688 454142
rect 517552 452460 518688 453604
rect 517552 451948 517606 452460
rect 518658 451948 518688 452460
rect 517552 451938 518688 451948
rect 522126 454970 522696 454978
rect 522126 454412 522198 454970
rect 522690 454412 522696 454970
rect 522126 450880 522696 454412
rect 522988 454970 523420 454976
rect 522988 454412 522994 454970
rect 523414 454412 523420 454970
rect 522988 454406 523420 454412
rect 522999 454142 523408 454154
rect 522999 453604 523005 454142
rect 523402 453604 523408 454142
rect 522999 453592 523408 453604
rect 522937 451688 523346 451700
rect 522937 451150 522943 451688
rect 523340 451150 523346 451688
rect 522937 451138 523346 451150
rect 522126 450322 522132 450880
rect 522690 450322 522696 450880
rect 522126 450316 522696 450322
rect 522926 450880 523358 450886
rect 522926 450322 522932 450880
rect 523352 450322 523358 450880
rect 522926 450316 523358 450322
rect 516852 448686 516858 449244
rect 517416 448686 517422 449244
rect 516852 448680 517422 448686
rect 517652 450062 518222 450068
rect 517652 449504 517658 450062
rect 518216 449504 518222 450062
rect 515390 447868 515396 448426
rect 515954 447868 515960 448426
rect 515390 447862 515960 447868
rect 516190 448426 516622 448432
rect 516190 447868 516196 448426
rect 516616 447868 516622 448426
rect 516190 447862 516622 447868
rect 514234 447616 514588 447816
rect 514788 447616 514926 447816
rect 514234 447416 514926 447616
rect 514234 447216 514588 447416
rect 514788 447216 514926 447416
rect 514234 447016 514926 447216
rect 516190 447608 516622 447614
rect 516190 447050 516196 447608
rect 516616 447050 516622 447608
rect 516190 447044 516622 447050
rect 516852 447608 517422 447614
rect 516852 447050 516858 447608
rect 517416 447050 517422 447608
rect 514234 446816 514588 447016
rect 514788 446816 514926 447016
rect 514234 446616 514926 446816
rect 514234 446416 514588 446616
rect 514788 446416 514926 446616
rect 503039 446308 503085 446320
rect 503039 446302 503045 446308
rect 502808 446282 503045 446302
rect 502808 446142 502828 446282
rect 502948 446142 503045 446282
rect 502808 446124 503045 446142
rect 503079 446302 503085 446308
rect 503079 446124 503088 446302
rect 502808 446122 503088 446124
rect 514234 446216 514926 446416
rect 516190 446790 516622 446796
rect 516190 446232 516196 446790
rect 516616 446232 516622 446790
rect 516190 446226 516622 446232
rect 503039 446112 503085 446122
rect 502648 446022 502768 446042
rect 502648 445942 502668 446022
rect 502748 446002 502768 446022
rect 514234 446016 514588 446216
rect 514788 446016 514926 446216
rect 503126 446004 510866 446010
rect 503126 446002 503138 446004
rect 502748 445970 503138 446002
rect 510854 445970 510866 446004
rect 502748 445964 510866 445970
rect 502748 445962 503148 445964
rect 502748 445942 502768 445962
rect 502648 445922 502768 445942
rect 503039 445850 503085 445862
rect 503039 445842 503045 445850
rect 502808 445822 503045 445842
rect 502808 445682 502828 445822
rect 502948 445682 503045 445822
rect 502808 445666 503045 445682
rect 503079 445842 503085 445850
rect 503079 445666 503088 445842
rect 502808 445662 503088 445666
rect 514234 445816 514926 446016
rect 503039 445654 503085 445662
rect 510928 445636 513328 445642
rect 510928 445562 512134 445636
rect 510828 445552 512134 445562
rect 503126 445546 512134 445552
rect 503126 445512 503138 445546
rect 510854 445512 512134 445546
rect 503126 445506 512134 445512
rect 510828 445502 512134 445506
rect 503039 445392 503085 445404
rect 503039 445382 503045 445392
rect 502808 445362 503045 445382
rect 502808 445222 502828 445362
rect 502948 445222 503045 445362
rect 502808 445208 503045 445222
rect 503079 445382 503085 445392
rect 503079 445208 503088 445382
rect 502808 445202 503088 445208
rect 503039 445196 503085 445202
rect 502648 445102 502768 445122
rect 502648 445022 502668 445102
rect 502748 445094 503148 445102
rect 502748 445088 510866 445094
rect 502748 445062 503138 445088
rect 502748 445022 502768 445062
rect 503126 445054 503138 445062
rect 510854 445054 510866 445088
rect 503126 445048 510866 445054
rect 502648 445002 502768 445022
rect 503039 444934 503085 444946
rect 503039 444922 503045 444934
rect 502808 444902 503045 444922
rect 502808 444762 502828 444902
rect 502948 444762 503045 444902
rect 502808 444750 503045 444762
rect 503079 444922 503085 444934
rect 503079 444750 503088 444922
rect 502808 444742 503088 444750
rect 503039 444738 503085 444742
rect 510928 444642 512134 445502
rect 510848 444636 512134 444642
rect 503126 444630 512134 444636
rect 503126 444596 503138 444630
rect 510854 444596 512134 444630
rect 503126 444590 512134 444596
rect 510848 444582 512134 444590
rect 503039 444476 503085 444488
rect 503039 444462 503045 444476
rect 502808 444442 503045 444462
rect 502808 444302 502828 444442
rect 502948 444302 503045 444442
rect 502808 444292 503045 444302
rect 503079 444462 503085 444476
rect 503079 444292 503088 444462
rect 502808 444282 503088 444292
rect 503039 444280 503085 444282
rect 502648 444182 502768 444202
rect 502648 444102 502668 444182
rect 502748 444178 503148 444182
rect 502748 444172 510866 444178
rect 502748 444142 503138 444172
rect 502748 444102 502768 444142
rect 503126 444138 503138 444142
rect 510854 444138 510866 444172
rect 503126 444132 510866 444138
rect 502648 444082 502768 444102
rect 503039 444018 503085 444030
rect 503039 444002 503045 444018
rect 502808 443982 503045 444002
rect 502808 443842 502828 443982
rect 502948 443842 503045 443982
rect 502808 443834 503045 443842
rect 503079 444002 503085 444018
rect 503079 443834 503088 444002
rect 502808 443822 503088 443834
rect 510928 443722 512134 444582
rect 510848 443720 512134 443722
rect 503122 443714 512134 443720
rect 503122 443680 503138 443714
rect 510854 443682 512134 443714
rect 510854 443680 510866 443682
rect 503122 443674 510866 443680
rect 502426 443560 503086 443674
rect 510928 443648 512134 443682
rect 512422 443648 512836 445636
rect 513286 443648 513328 445636
rect 510928 443642 513328 443648
rect 514234 445616 514588 445816
rect 514788 445616 514926 445816
rect 514234 444216 514926 445616
rect 514234 444016 514588 444216
rect 514788 444016 514926 444216
rect 514234 443816 514926 444016
rect 502426 443376 503045 443560
rect 503079 443376 503086 443560
rect 502426 443262 503086 443376
rect 514234 443616 514588 443816
rect 514788 443616 514926 443816
rect 514234 443416 514926 443616
rect 502426 443256 510866 443262
rect 502426 443222 503138 443256
rect 510854 443222 510866 443256
rect 502426 443216 510866 443222
rect 514234 443216 514588 443416
rect 514788 443216 514926 443416
rect 502426 442986 502726 443216
rect 502426 442586 502526 442986
rect 502626 442586 502726 442986
rect 502426 442486 502726 442586
rect 514234 443016 514926 443216
rect 514234 442816 514588 443016
rect 514788 442816 514926 443016
rect 514234 442616 514926 442816
rect 514234 442416 514588 442616
rect 514788 442416 514926 442616
rect 514234 442216 514926 442416
rect 514234 442016 514588 442216
rect 514788 442016 514926 442216
rect 515390 445972 515960 445978
rect 515390 445414 515396 445972
rect 515954 445414 515960 445972
rect 515390 442700 515960 445414
rect 516190 445972 516622 445978
rect 516190 445414 516196 445972
rect 516616 445414 516622 445972
rect 516190 445408 516622 445414
rect 516066 445232 516622 445238
rect 516584 445154 516622 445232
rect 516616 444596 516622 445154
rect 516584 444540 516622 444596
rect 516066 444534 516622 444540
rect 516190 444336 516622 444342
rect 516190 443778 516196 444336
rect 516616 443778 516622 444336
rect 516190 443772 516622 443778
rect 516190 443518 516622 443524
rect 516190 442960 516196 443518
rect 516616 442960 516622 443518
rect 516190 442954 516622 442960
rect 516852 443518 517422 447050
rect 517652 446790 518222 449504
rect 522926 450062 523358 450068
rect 522926 449504 522932 450062
rect 523352 449504 523358 450062
rect 522926 449498 523358 449504
rect 523588 450062 524158 455230
rect 562150 455440 567584 455473
rect 562150 455360 562480 455440
rect 562560 455360 562640 455440
rect 562720 455360 562800 455440
rect 562880 455360 562960 455440
rect 563040 455360 563120 455440
rect 563200 455360 563280 455440
rect 563360 455360 563440 455440
rect 563520 455360 563600 455440
rect 563680 455360 563760 455440
rect 563840 455360 563920 455440
rect 564000 455360 564080 455440
rect 564160 455360 564240 455440
rect 564320 455360 564400 455440
rect 564480 455360 564560 455440
rect 564640 455360 564720 455440
rect 564800 455360 564880 455440
rect 564960 455360 565040 455440
rect 565120 455360 565200 455440
rect 565280 455360 565360 455440
rect 565440 455360 565520 455440
rect 565600 455360 565680 455440
rect 565760 455360 565840 455440
rect 565920 455360 566000 455440
rect 566080 455360 566160 455440
rect 566240 455360 566320 455440
rect 566400 455360 566480 455440
rect 566560 455360 566640 455440
rect 566720 455360 566800 455440
rect 566880 455360 566960 455440
rect 567040 455360 567120 455440
rect 567200 455360 567280 455440
rect 567360 455360 567584 455440
rect 562150 455280 567584 455360
rect 562150 455212 562480 455280
rect 562560 455212 562640 455280
rect 562720 455212 562800 455280
rect 562880 455212 562960 455280
rect 563040 455212 563120 455280
rect 563200 455212 563280 455280
rect 563360 455212 563440 455280
rect 563520 455212 563600 455280
rect 563680 455212 563760 455280
rect 563840 455212 563920 455280
rect 564000 455212 564080 455280
rect 564160 455212 564240 455280
rect 564320 455212 564400 455280
rect 564480 455212 564560 455280
rect 564640 455212 564720 455280
rect 564800 455212 564880 455280
rect 564960 455212 565040 455280
rect 565120 455212 565200 455280
rect 565280 455212 565360 455280
rect 565440 455212 565520 455280
rect 565600 455212 565680 455280
rect 565760 455212 565840 455280
rect 565920 455212 566000 455280
rect 566080 455212 566160 455280
rect 566240 455212 566320 455280
rect 566400 455212 566480 455280
rect 566560 455212 566640 455280
rect 566720 455212 566800 455280
rect 566880 455212 566960 455280
rect 567040 455212 567120 455280
rect 567200 455212 567280 455280
rect 567360 455212 567584 455280
rect 562150 455178 562190 455212
rect 567544 455178 567584 455212
rect 562150 455172 567584 455178
rect 562150 455055 562196 455172
rect 562150 454073 562156 455055
rect 562190 454073 562196 455055
rect 562150 454061 562196 454073
rect 562264 455088 562310 455100
rect 562264 454112 562270 455088
rect 562304 454112 562310 455088
rect 562264 453975 562310 454112
rect 562522 455088 562568 455172
rect 562522 454112 562528 455088
rect 562562 454112 562568 455088
rect 562522 454100 562568 454112
rect 562780 455088 562826 455100
rect 562780 454112 562786 455088
rect 562820 454112 562826 455088
rect 562362 454053 562470 454059
rect 562362 454019 562374 454053
rect 562458 454019 562470 454053
rect 562362 454013 562470 454019
rect 562620 454053 562728 454059
rect 562620 454019 562632 454053
rect 562716 454019 562728 454053
rect 562620 454013 562728 454019
rect 562780 453975 562826 454112
rect 563038 455088 563084 455172
rect 563038 454112 563044 455088
rect 563078 454112 563084 455088
rect 563038 454100 563084 454112
rect 563296 455088 563342 455100
rect 563296 454112 563302 455088
rect 563336 454112 563342 455088
rect 562878 454053 562986 454059
rect 562878 454019 562890 454053
rect 562974 454019 562986 454053
rect 562878 454013 562986 454019
rect 563136 454053 563244 454059
rect 563136 454019 563148 454053
rect 563232 454019 563244 454053
rect 563136 454013 563244 454019
rect 563296 453975 563342 454112
rect 563554 455088 563600 455172
rect 563554 454112 563560 455088
rect 563594 454112 563600 455088
rect 563554 454100 563600 454112
rect 563812 455088 563858 455100
rect 563812 454112 563818 455088
rect 563852 454112 563858 455088
rect 563394 454053 563502 454059
rect 563394 454019 563406 454053
rect 563490 454019 563502 454053
rect 563394 454013 563502 454019
rect 563652 454053 563760 454059
rect 563652 454019 563664 454053
rect 563748 454019 563760 454053
rect 563652 454013 563760 454019
rect 563812 453975 563858 454112
rect 564070 455088 564116 455172
rect 564070 454112 564076 455088
rect 564110 454112 564116 455088
rect 564070 454100 564116 454112
rect 564328 455088 564374 455100
rect 564328 454112 564334 455088
rect 564368 454112 564374 455088
rect 563910 454053 564018 454059
rect 563910 454019 563922 454053
rect 564006 454019 564018 454053
rect 563910 454013 564018 454019
rect 564168 454053 564276 454059
rect 564168 454019 564180 454053
rect 564264 454019 564276 454053
rect 564168 454013 564276 454019
rect 564328 453975 564374 454112
rect 564586 455088 564632 455172
rect 564586 454112 564592 455088
rect 564626 454112 564632 455088
rect 564586 454100 564632 454112
rect 564844 455088 564890 455100
rect 564844 454112 564850 455088
rect 564884 454112 564890 455088
rect 564426 454053 564534 454059
rect 564426 454019 564438 454053
rect 564522 454019 564534 454053
rect 564426 454013 564534 454019
rect 564684 454053 564792 454059
rect 564684 454019 564696 454053
rect 564780 454019 564792 454053
rect 564684 454013 564792 454019
rect 564844 453975 564890 454112
rect 565102 455088 565148 455172
rect 565102 454112 565108 455088
rect 565142 454112 565148 455088
rect 565102 454100 565148 454112
rect 565360 455088 565406 455100
rect 565360 454112 565366 455088
rect 565400 454112 565406 455088
rect 564942 454053 565050 454059
rect 564942 454019 564954 454053
rect 565038 454019 565050 454053
rect 564942 454013 565050 454019
rect 565200 454053 565308 454059
rect 565200 454019 565212 454053
rect 565296 454019 565308 454053
rect 565200 454013 565308 454019
rect 565360 453975 565406 454112
rect 565618 455088 565664 455172
rect 565618 454112 565624 455088
rect 565658 454112 565664 455088
rect 565618 454100 565664 454112
rect 565876 455088 565922 455100
rect 565876 454112 565882 455088
rect 565916 454112 565922 455088
rect 565458 454053 565566 454059
rect 565458 454019 565470 454053
rect 565554 454019 565566 454053
rect 565458 454013 565566 454019
rect 565716 454053 565824 454059
rect 565716 454019 565728 454053
rect 565812 454019 565824 454053
rect 565716 454013 565824 454019
rect 565876 453975 565922 454112
rect 566134 455088 566180 455172
rect 566134 454112 566140 455088
rect 566174 454112 566180 455088
rect 566134 454100 566180 454112
rect 566392 455088 566438 455100
rect 566392 454112 566398 455088
rect 566432 454112 566438 455088
rect 565974 454053 566082 454059
rect 565974 454019 565986 454053
rect 566070 454019 566082 454053
rect 565974 454013 566082 454019
rect 566232 454053 566340 454059
rect 566232 454019 566244 454053
rect 566328 454019 566340 454053
rect 566232 454013 566340 454019
rect 566392 453975 566438 454112
rect 566650 455088 566696 455172
rect 566650 454112 566656 455088
rect 566690 454112 566696 455088
rect 566650 454100 566696 454112
rect 566908 455088 566954 455100
rect 566908 454112 566914 455088
rect 566948 454112 566954 455088
rect 566490 454053 566598 454059
rect 566490 454019 566502 454053
rect 566586 454019 566598 454053
rect 566490 454013 566598 454019
rect 566748 454053 566856 454059
rect 566748 454019 566760 454053
rect 566844 454019 566856 454053
rect 566748 454013 566856 454019
rect 566908 453975 566954 454112
rect 567166 455088 567212 455172
rect 567166 454112 567172 455088
rect 567206 454112 567212 455088
rect 567166 454100 567212 454112
rect 567424 455088 567470 455100
rect 567424 454112 567430 455088
rect 567464 454112 567470 455088
rect 567006 454053 567114 454059
rect 567006 454019 567018 454053
rect 567102 454019 567114 454053
rect 567006 454013 567114 454019
rect 567264 454053 567372 454059
rect 567264 454019 567276 454053
rect 567360 454019 567372 454053
rect 567264 454013 567372 454019
rect 567424 453975 567470 454112
rect 567538 455055 567584 455172
rect 567538 454073 567544 455055
rect 567578 454073 567584 455055
rect 572310 455440 577744 455473
rect 572310 455360 572640 455440
rect 572720 455360 572800 455440
rect 572880 455360 572960 455440
rect 573040 455360 573120 455440
rect 573200 455360 573280 455440
rect 573360 455360 573440 455440
rect 573520 455360 573600 455440
rect 573680 455360 573760 455440
rect 573840 455360 573920 455440
rect 574000 455360 574080 455440
rect 574160 455360 574240 455440
rect 574320 455360 574400 455440
rect 574480 455360 574560 455440
rect 574640 455360 574720 455440
rect 574800 455360 574880 455440
rect 574960 455360 575040 455440
rect 575120 455360 575200 455440
rect 575280 455360 575360 455440
rect 575440 455360 575520 455440
rect 575600 455360 575680 455440
rect 575760 455360 575840 455440
rect 575920 455360 576000 455440
rect 576080 455360 576160 455440
rect 576240 455360 576320 455440
rect 576400 455360 576480 455440
rect 576560 455360 576640 455440
rect 576720 455360 576800 455440
rect 576880 455360 576960 455440
rect 577040 455360 577120 455440
rect 577200 455360 577280 455440
rect 577360 455360 577440 455440
rect 577520 455360 577744 455440
rect 572310 455280 577744 455360
rect 572310 455246 572640 455280
rect 572720 455246 572800 455280
rect 572880 455246 572960 455280
rect 573040 455246 573120 455280
rect 573200 455246 573280 455280
rect 573360 455246 573440 455280
rect 573520 455246 573600 455280
rect 573680 455246 573760 455280
rect 573840 455246 573920 455280
rect 574000 455246 574080 455280
rect 574160 455246 574240 455280
rect 574320 455246 574400 455280
rect 574480 455246 574560 455280
rect 574640 455246 574720 455280
rect 574800 455246 574880 455280
rect 574960 455246 575040 455280
rect 575120 455246 575200 455280
rect 575280 455246 575360 455280
rect 575440 455246 575520 455280
rect 575600 455246 575680 455280
rect 575760 455246 575840 455280
rect 575920 455246 576000 455280
rect 576080 455246 576160 455280
rect 576240 455246 576320 455280
rect 576400 455246 576480 455280
rect 576560 455246 576640 455280
rect 576720 455246 576800 455280
rect 576880 455246 576960 455280
rect 577040 455246 577120 455280
rect 577200 455246 577280 455280
rect 577360 455246 577440 455280
rect 577520 455246 577744 455280
rect 572310 455212 572350 455246
rect 577704 455212 577744 455246
rect 572310 455200 572640 455212
rect 572720 455200 572800 455212
rect 572880 455200 572960 455212
rect 573040 455200 573120 455212
rect 573200 455200 573280 455212
rect 573360 455200 573440 455212
rect 573520 455200 573600 455212
rect 573680 455200 573760 455212
rect 573840 455200 573920 455212
rect 574000 455200 574080 455212
rect 574160 455200 574240 455212
rect 574320 455200 574400 455212
rect 574480 455200 574560 455212
rect 574640 455200 574720 455212
rect 574800 455200 574880 455212
rect 574960 455200 575040 455212
rect 575120 455200 575200 455212
rect 575280 455200 575360 455212
rect 575440 455200 575520 455212
rect 575600 455200 575680 455212
rect 575760 455200 575840 455212
rect 575920 455200 576000 455212
rect 576080 455200 576160 455212
rect 576240 455200 576320 455212
rect 576400 455200 576480 455212
rect 576560 455200 576640 455212
rect 576720 455200 576800 455212
rect 576880 455200 576960 455212
rect 577040 455200 577120 455212
rect 577200 455200 577280 455212
rect 577360 455200 577440 455212
rect 577520 455200 577744 455212
rect 572310 455172 577744 455200
rect 572310 455090 572356 455172
rect 572688 455134 572722 455172
rect 573204 455134 573238 455172
rect 573720 455134 573754 455172
rect 574236 455134 574270 455172
rect 574752 455134 574786 455172
rect 575268 455134 575302 455172
rect 575784 455134 575818 455172
rect 576300 455134 576334 455172
rect 576816 455134 576850 455172
rect 577332 455134 577366 455172
rect 572310 454116 572316 455090
rect 572350 454116 572356 455090
rect 572310 454104 572356 454116
rect 572424 455122 572470 455134
rect 572424 454146 572430 455122
rect 572464 454146 572470 455122
rect 567538 454061 567584 454073
rect 572424 453990 572470 454146
rect 572682 455122 572728 455134
rect 572682 454146 572688 455122
rect 572722 454146 572728 455122
rect 572682 454134 572728 454146
rect 572940 455122 572986 455134
rect 572940 454146 572946 455122
rect 572980 454146 572986 455122
rect 572522 454096 572630 454102
rect 572522 454062 572534 454096
rect 572618 454062 572630 454096
rect 572522 454056 572630 454062
rect 572780 454096 572888 454102
rect 572780 454062 572792 454096
rect 572876 454062 572888 454096
rect 572780 454056 572888 454062
rect 572940 453990 572986 454146
rect 573198 455122 573244 455134
rect 573198 454146 573204 455122
rect 573238 454146 573244 455122
rect 573198 454134 573244 454146
rect 573456 455122 573502 455134
rect 573456 454146 573462 455122
rect 573496 454146 573502 455122
rect 573038 454096 573146 454102
rect 573038 454062 573050 454096
rect 573134 454062 573146 454096
rect 573038 454056 573146 454062
rect 573296 454096 573404 454102
rect 573296 454062 573308 454096
rect 573392 454062 573404 454096
rect 573296 454056 573404 454062
rect 573456 453990 573502 454146
rect 573714 455122 573760 455134
rect 573714 454146 573720 455122
rect 573754 454146 573760 455122
rect 573714 454134 573760 454146
rect 573972 455122 574018 455134
rect 573972 454146 573978 455122
rect 574012 454146 574018 455122
rect 573554 454096 573662 454102
rect 573554 454062 573566 454096
rect 573650 454062 573662 454096
rect 573554 454056 573662 454062
rect 573812 454096 573920 454102
rect 573812 454062 573824 454096
rect 573908 454062 573920 454096
rect 573812 454056 573920 454062
rect 573972 453990 574018 454146
rect 574230 455122 574276 455134
rect 574230 454146 574236 455122
rect 574270 454146 574276 455122
rect 574230 454134 574276 454146
rect 574488 455122 574534 455134
rect 574488 454146 574494 455122
rect 574528 454146 574534 455122
rect 574070 454096 574178 454102
rect 574070 454062 574082 454096
rect 574166 454062 574178 454096
rect 574070 454056 574178 454062
rect 574328 454096 574436 454102
rect 574328 454062 574340 454096
rect 574424 454062 574436 454096
rect 574328 454056 574436 454062
rect 574488 453990 574534 454146
rect 574746 455122 574792 455134
rect 574746 454146 574752 455122
rect 574786 454146 574792 455122
rect 574746 454134 574792 454146
rect 575004 455122 575050 455134
rect 575004 454146 575010 455122
rect 575044 454146 575050 455122
rect 574586 454096 574694 454102
rect 574586 454062 574598 454096
rect 574682 454062 574694 454096
rect 574586 454056 574694 454062
rect 574844 454096 574952 454102
rect 574844 454062 574856 454096
rect 574940 454062 574952 454096
rect 574844 454056 574952 454062
rect 575004 453990 575050 454146
rect 575262 455122 575308 455134
rect 575262 454146 575268 455122
rect 575302 454146 575308 455122
rect 575262 454134 575308 454146
rect 575520 455122 575566 455134
rect 575520 454146 575526 455122
rect 575560 454146 575566 455122
rect 575102 454096 575210 454102
rect 575102 454062 575114 454096
rect 575198 454062 575210 454096
rect 575102 454056 575210 454062
rect 575360 454096 575468 454102
rect 575360 454062 575372 454096
rect 575456 454062 575468 454096
rect 575360 454056 575468 454062
rect 575520 453990 575566 454146
rect 575778 455122 575824 455134
rect 575778 454146 575784 455122
rect 575818 454146 575824 455122
rect 575778 454134 575824 454146
rect 576036 455122 576082 455134
rect 576036 454146 576042 455122
rect 576076 454146 576082 455122
rect 575618 454096 575726 454102
rect 575618 454062 575630 454096
rect 575714 454062 575726 454096
rect 575618 454056 575726 454062
rect 575876 454096 575984 454102
rect 575876 454062 575888 454096
rect 575972 454062 575984 454096
rect 575876 454056 575984 454062
rect 576036 453990 576082 454146
rect 576294 455122 576340 455134
rect 576294 454146 576300 455122
rect 576334 454146 576340 455122
rect 576294 454134 576340 454146
rect 576552 455122 576598 455134
rect 576552 454146 576558 455122
rect 576592 454146 576598 455122
rect 576134 454096 576242 454102
rect 576134 454062 576146 454096
rect 576230 454062 576242 454096
rect 576134 454056 576242 454062
rect 576392 454096 576500 454102
rect 576392 454062 576404 454096
rect 576488 454062 576500 454096
rect 576392 454056 576500 454062
rect 576552 453990 576598 454146
rect 576810 455122 576856 455134
rect 576810 454146 576816 455122
rect 576850 454146 576856 455122
rect 576810 454134 576856 454146
rect 577068 455122 577114 455134
rect 577068 454146 577074 455122
rect 577108 454146 577114 455122
rect 576650 454096 576758 454102
rect 576650 454062 576662 454096
rect 576746 454062 576758 454096
rect 576650 454056 576758 454062
rect 576908 454096 577016 454102
rect 576908 454062 576920 454096
rect 577004 454062 577016 454096
rect 576908 454056 577016 454062
rect 577068 453990 577114 454146
rect 577326 455122 577372 455134
rect 577326 454146 577332 455122
rect 577366 454146 577372 455122
rect 577326 454134 577372 454146
rect 577584 455122 577630 455134
rect 577584 454146 577590 455122
rect 577624 454146 577630 455122
rect 577166 454096 577274 454102
rect 577166 454062 577178 454096
rect 577262 454062 577274 454096
rect 577166 454056 577274 454062
rect 577424 454096 577532 454102
rect 577424 454062 577436 454096
rect 577520 454062 577532 454096
rect 577424 454056 577532 454062
rect 577584 453990 577630 454146
rect 577698 455090 577744 455172
rect 577698 454116 577704 455090
rect 577738 454116 577744 455090
rect 577698 454104 577744 454116
rect 562120 453919 567614 453975
rect 562120 453859 562222 453919
rect 562282 453859 562342 453919
rect 562402 453859 562462 453919
rect 562522 453859 562582 453919
rect 562642 453859 562702 453919
rect 562762 453859 562822 453919
rect 562882 453859 562942 453919
rect 563002 453859 563062 453919
rect 563122 453859 563182 453919
rect 563242 453859 563302 453919
rect 563362 453859 563422 453919
rect 563482 453859 563542 453919
rect 563602 453859 563662 453919
rect 563722 453859 563782 453919
rect 563842 453859 563902 453919
rect 563962 453859 564022 453919
rect 564082 453859 564142 453919
rect 564202 453859 564262 453919
rect 564322 453859 564382 453919
rect 564442 453859 564502 453919
rect 564562 453859 564622 453919
rect 564682 453859 564742 453919
rect 564802 453859 564862 453919
rect 564922 453859 564982 453919
rect 565042 453859 565102 453919
rect 565162 453859 565222 453919
rect 565282 453859 565342 453919
rect 565402 453859 565462 453919
rect 565522 453859 565582 453919
rect 565642 453859 565702 453919
rect 565762 453859 565822 453919
rect 565882 453859 565942 453919
rect 566002 453859 566062 453919
rect 566122 453859 566182 453919
rect 566242 453859 566302 453919
rect 566362 453859 566422 453919
rect 566482 453859 566542 453919
rect 566602 453859 566662 453919
rect 566722 453859 566782 453919
rect 566842 453859 566902 453919
rect 566962 453859 567022 453919
rect 567082 453859 567142 453919
rect 567202 453859 567262 453919
rect 567322 453859 567382 453919
rect 567442 453859 567502 453919
rect 567562 453859 567614 453919
rect 562120 453799 567614 453859
rect 562120 453739 562222 453799
rect 562282 453739 562342 453799
rect 562402 453739 562462 453799
rect 562522 453739 562582 453799
rect 562642 453739 562702 453799
rect 562762 453739 562822 453799
rect 562882 453739 562942 453799
rect 563002 453739 563062 453799
rect 563122 453739 563182 453799
rect 563242 453739 563302 453799
rect 563362 453739 563422 453799
rect 563482 453739 563542 453799
rect 563602 453739 563662 453799
rect 563722 453739 563782 453799
rect 563842 453739 563902 453799
rect 563962 453739 564022 453799
rect 564082 453739 564142 453799
rect 564202 453739 564262 453799
rect 564322 453739 564382 453799
rect 564442 453739 564502 453799
rect 564562 453739 564622 453799
rect 564682 453739 564742 453799
rect 564802 453739 564862 453799
rect 564922 453739 564982 453799
rect 565042 453739 565102 453799
rect 565162 453739 565222 453799
rect 565282 453739 565342 453799
rect 565402 453739 565462 453799
rect 565522 453739 565582 453799
rect 565642 453739 565702 453799
rect 565762 453739 565822 453799
rect 565882 453739 565942 453799
rect 566002 453739 566062 453799
rect 566122 453739 566182 453799
rect 566242 453739 566302 453799
rect 566362 453739 566422 453799
rect 566482 453739 566542 453799
rect 566602 453739 566662 453799
rect 566722 453739 566782 453799
rect 566842 453739 566902 453799
rect 566962 453739 567022 453799
rect 567082 453739 567142 453799
rect 567202 453739 567262 453799
rect 567322 453739 567382 453799
rect 567442 453739 567502 453799
rect 567562 453739 567614 453799
rect 562120 453700 567614 453739
rect 572280 453934 577774 453990
rect 572280 453874 572332 453934
rect 572392 453874 572452 453934
rect 572512 453874 572572 453934
rect 572632 453874 572692 453934
rect 572752 453874 572812 453934
rect 572872 453874 572932 453934
rect 572992 453874 573052 453934
rect 573112 453874 573172 453934
rect 573232 453874 573292 453934
rect 573352 453874 573412 453934
rect 573472 453874 573532 453934
rect 573592 453874 573652 453934
rect 573712 453874 573772 453934
rect 573832 453874 573892 453934
rect 573952 453874 574012 453934
rect 574072 453874 574132 453934
rect 574192 453874 574252 453934
rect 574312 453874 574372 453934
rect 574432 453874 574492 453934
rect 574552 453874 574612 453934
rect 574672 453874 574732 453934
rect 574792 453874 574852 453934
rect 574912 453874 574972 453934
rect 575032 453874 575092 453934
rect 575152 453874 575212 453934
rect 575272 453874 575332 453934
rect 575392 453874 575452 453934
rect 575512 453874 575572 453934
rect 575632 453874 575692 453934
rect 575752 453874 575812 453934
rect 575872 453874 575932 453934
rect 575992 453874 576052 453934
rect 576112 453874 576172 453934
rect 576232 453874 576292 453934
rect 576352 453874 576412 453934
rect 576472 453874 576532 453934
rect 576592 453874 576652 453934
rect 576712 453874 576772 453934
rect 576832 453874 576892 453934
rect 576952 453874 577012 453934
rect 577072 453874 577132 453934
rect 577192 453874 577252 453934
rect 577312 453874 577372 453934
rect 577432 453874 577492 453934
rect 577552 453874 577612 453934
rect 577672 453874 577774 453934
rect 572280 453814 577774 453874
rect 572280 453754 572332 453814
rect 572392 453754 572452 453814
rect 572512 453754 572572 453814
rect 572632 453754 572692 453814
rect 572752 453754 572812 453814
rect 572872 453754 572932 453814
rect 572992 453754 573052 453814
rect 573112 453754 573172 453814
rect 573232 453754 573292 453814
rect 573352 453754 573412 453814
rect 573472 453754 573532 453814
rect 573592 453754 573652 453814
rect 573712 453754 573772 453814
rect 573832 453754 573892 453814
rect 573952 453754 574012 453814
rect 574072 453754 574132 453814
rect 574192 453754 574252 453814
rect 574312 453754 574372 453814
rect 574432 453754 574492 453814
rect 574552 453754 574612 453814
rect 574672 453754 574732 453814
rect 574792 453754 574852 453814
rect 574912 453754 574972 453814
rect 575032 453754 575092 453814
rect 575152 453754 575212 453814
rect 575272 453754 575332 453814
rect 575392 453754 575452 453814
rect 575512 453754 575572 453814
rect 575632 453754 575692 453814
rect 575752 453754 575812 453814
rect 575872 453754 575932 453814
rect 575992 453754 576052 453814
rect 576112 453754 576172 453814
rect 576232 453754 576292 453814
rect 576352 453754 576412 453814
rect 576472 453754 576532 453814
rect 576592 453754 576652 453814
rect 576712 453754 576772 453814
rect 576832 453754 576892 453814
rect 576952 453754 577012 453814
rect 577072 453754 577132 453814
rect 577192 453754 577252 453814
rect 577312 453754 577372 453814
rect 577432 453754 577492 453814
rect 577552 453754 577612 453814
rect 577672 453754 577774 453814
rect 572280 453715 577774 453754
rect 523588 449504 523594 450062
rect 524152 449504 524158 450062
rect 523588 449498 524158 449504
rect 522926 449244 523358 449250
rect 522926 448686 522932 449244
rect 523352 448686 523358 449244
rect 522926 448680 523358 448686
rect 524388 449232 524958 449238
rect 524388 448674 524394 449232
rect 524952 448674 524958 449232
rect 517652 446232 517658 446790
rect 518216 446232 518222 446790
rect 517652 446226 518222 446232
rect 522126 448426 522696 448432
rect 522126 447868 522132 448426
rect 522690 447868 522696 448426
rect 522126 445972 522696 447868
rect 522926 448426 523358 448432
rect 522926 447868 522932 448426
rect 523352 447868 523358 448426
rect 522926 447862 523358 447868
rect 522926 447608 523358 447614
rect 522926 447050 522932 447608
rect 523352 447050 523358 447608
rect 522926 447044 523358 447050
rect 524388 447608 524958 448674
rect 524388 447050 524394 447608
rect 524952 447050 524958 447608
rect 524388 447044 524958 447050
rect 522926 446790 523358 446796
rect 522926 446232 522932 446790
rect 523352 446232 523358 446790
rect 522926 446226 523358 446232
rect 523588 446790 524158 446918
rect 523588 446232 523594 446790
rect 524152 446232 524158 446790
rect 522126 445414 522132 445972
rect 522690 445414 522696 445972
rect 522126 445408 522696 445414
rect 522926 445972 523358 445978
rect 522926 445414 522932 445972
rect 523352 445414 523358 445972
rect 522926 445408 523358 445414
rect 522926 445154 523358 445160
rect 522926 444596 522932 445154
rect 523352 444596 523358 445154
rect 522926 444590 523358 444596
rect 522926 444336 523358 444342
rect 516852 442960 516858 443518
rect 517416 442960 517422 443518
rect 516852 442954 517422 442960
rect 517652 443778 517658 444336
rect 518216 443778 518222 444336
rect 515390 442142 515396 442700
rect 515954 442142 515960 442700
rect 515390 442136 515960 442142
rect 516190 442700 516622 442706
rect 516190 442142 516196 442700
rect 516616 442142 516622 442700
rect 516190 442136 516622 442142
rect 514234 441816 514926 442016
rect 503646 441668 514072 441674
rect 503646 440732 503652 441668
rect 504588 441666 514072 441668
rect 504588 440732 513548 441666
rect 514066 440732 514072 441666
rect 503646 440726 514072 440732
rect 514234 441616 514588 441816
rect 514788 441616 514926 441816
rect 514234 441416 514926 441616
rect 514234 441216 514588 441416
rect 514788 441216 514926 441416
rect 516190 441882 516622 441888
rect 516190 441324 516196 441882
rect 516616 441324 516622 441882
rect 516190 441318 516622 441324
rect 517652 441882 518222 443778
rect 522926 443778 522932 444336
rect 523352 443778 523358 444336
rect 522926 443772 523358 443778
rect 523588 444336 524158 446232
rect 523588 443778 523594 444336
rect 524152 443778 524158 444336
rect 523588 443772 524158 443778
rect 522926 443518 523358 443524
rect 522926 442960 522932 443518
rect 523352 442960 523358 443518
rect 522926 442954 523358 442960
rect 524388 443518 524958 443692
rect 524388 442960 524394 443518
rect 524952 442960 524958 443518
rect 517652 441324 517658 441882
rect 518216 441324 518222 441882
rect 517652 441318 518222 441324
rect 522126 442700 522696 442706
rect 522126 442142 522132 442700
rect 522690 442142 522696 442700
rect 514234 441148 514926 441216
rect 514234 441142 516622 441148
rect 514234 441016 515924 441142
rect 514234 440816 514588 441016
rect 514788 440816 515924 441016
rect 514234 440450 515924 440816
rect 516616 440450 516622 441142
rect 514234 440444 516622 440450
rect 508798 440324 516622 440330
rect 508798 439632 508806 440324
rect 509498 439632 512836 440324
rect 513286 439632 515924 440324
rect 516616 439632 516622 440324
rect 522126 440246 522696 442142
rect 522926 442700 523358 442706
rect 522926 442142 522932 442700
rect 523352 442142 523358 442700
rect 522926 442136 523358 442142
rect 522926 441882 523358 441888
rect 522926 441324 522932 441882
rect 523352 441324 523358 441882
rect 522926 441318 523358 441324
rect 523588 441882 524158 442002
rect 523588 441324 523594 441882
rect 524152 441324 524158 441882
rect 522926 441064 523358 441070
rect 522926 440506 522932 441064
rect 523352 440506 523358 441064
rect 522926 440500 523358 440506
rect 522126 439688 522132 440246
rect 522690 439688 522696 440246
rect 522126 439682 522696 439688
rect 522926 440246 523358 440252
rect 522926 439688 522932 440246
rect 523352 439688 523358 440246
rect 522926 439682 523358 439688
rect 508798 439626 516622 439632
rect 511528 439506 516622 439512
rect 511528 439504 515924 439506
rect 511528 438814 511534 439504
rect 511822 438814 515924 439504
rect 516616 438814 516622 439506
rect 522926 439428 523358 439434
rect 522926 438870 522932 439428
rect 523352 438870 523358 439428
rect 522926 438864 523358 438870
rect 523588 439428 524158 441324
rect 524388 441064 524958 442960
rect 524388 440506 524394 441064
rect 524952 440506 524958 441064
rect 524388 440494 524958 440506
rect 523588 438870 523594 439428
rect 524152 438870 524158 439428
rect 523588 438864 524158 438870
rect 511528 438808 516622 438814
rect 516202 438600 516611 438612
rect 503709 438112 513335 438143
rect 503709 438078 503740 438112
rect 503774 438078 503840 438112
rect 503874 438078 503940 438112
rect 503974 438078 504040 438112
rect 504074 438078 504140 438112
rect 504174 438078 504240 438112
rect 504274 438078 505028 438112
rect 505062 438078 505128 438112
rect 505162 438078 505228 438112
rect 505262 438078 505328 438112
rect 505362 438078 505428 438112
rect 505462 438078 505528 438112
rect 505562 438078 506316 438112
rect 506350 438078 506416 438112
rect 506450 438078 506516 438112
rect 506550 438078 506616 438112
rect 506650 438078 506716 438112
rect 506750 438078 506816 438112
rect 506850 438078 507604 438112
rect 507638 438078 507704 438112
rect 507738 438078 507804 438112
rect 507838 438078 507904 438112
rect 507938 438078 508004 438112
rect 508038 438078 508104 438112
rect 508138 438078 508892 438112
rect 508926 438078 508992 438112
rect 509026 438078 509092 438112
rect 509126 438078 509192 438112
rect 509226 438078 509292 438112
rect 509326 438078 509392 438112
rect 509426 438078 510180 438112
rect 510214 438078 510280 438112
rect 510314 438078 510380 438112
rect 510414 438078 510480 438112
rect 510514 438078 510580 438112
rect 510614 438078 510680 438112
rect 510714 438078 511468 438112
rect 511502 438078 511568 438112
rect 511602 438078 511668 438112
rect 511702 438078 511768 438112
rect 511802 438078 511868 438112
rect 511902 438078 511968 438112
rect 512002 438078 512756 438112
rect 512790 438078 512856 438112
rect 512890 438078 512956 438112
rect 512990 438078 513056 438112
rect 513090 438078 513156 438112
rect 513190 438078 513256 438112
rect 513290 438078 513335 438112
rect 503709 438012 513335 438078
rect 516202 438062 516208 438600
rect 516605 438062 516611 438600
rect 516202 438050 516611 438062
rect 522937 438600 523346 438612
rect 522937 438062 522943 438600
rect 523340 438062 523346 438600
rect 522937 438050 523346 438062
rect 503709 437978 503740 438012
rect 503774 437978 503840 438012
rect 503874 437978 503940 438012
rect 503974 437978 504040 438012
rect 504074 437978 504140 438012
rect 504174 437978 504240 438012
rect 504274 437978 505028 438012
rect 505062 437978 505128 438012
rect 505162 437978 505228 438012
rect 505262 437978 505328 438012
rect 505362 437978 505428 438012
rect 505462 437978 505528 438012
rect 505562 437978 506316 438012
rect 506350 437978 506416 438012
rect 506450 437978 506516 438012
rect 506550 437978 506616 438012
rect 506650 437978 506716 438012
rect 506750 437978 506816 438012
rect 506850 437978 507604 438012
rect 507638 437978 507704 438012
rect 507738 437978 507804 438012
rect 507838 437978 507904 438012
rect 507938 437978 508004 438012
rect 508038 437978 508104 438012
rect 508138 437978 508892 438012
rect 508926 437978 508992 438012
rect 509026 437978 509092 438012
rect 509126 437978 509192 438012
rect 509226 437978 509292 438012
rect 509326 437978 509392 438012
rect 509426 437978 510180 438012
rect 510214 437978 510280 438012
rect 510314 437978 510380 438012
rect 510414 437978 510480 438012
rect 510514 437978 510580 438012
rect 510614 437978 510680 438012
rect 510714 437978 511468 438012
rect 511502 437978 511568 438012
rect 511602 437978 511668 438012
rect 511702 437978 511768 438012
rect 511802 437978 511868 438012
rect 511902 437978 511968 438012
rect 512002 437978 512756 438012
rect 512790 437978 512856 438012
rect 512890 437978 512956 438012
rect 512990 437978 513056 438012
rect 513090 437978 513156 438012
rect 513190 437978 513256 438012
rect 513290 437978 513335 438012
rect 503709 437912 513335 437978
rect 503709 437878 503740 437912
rect 503774 437878 503840 437912
rect 503874 437878 503940 437912
rect 503974 437878 504040 437912
rect 504074 437878 504140 437912
rect 504174 437878 504240 437912
rect 504274 437878 505028 437912
rect 505062 437878 505128 437912
rect 505162 437878 505228 437912
rect 505262 437878 505328 437912
rect 505362 437878 505428 437912
rect 505462 437878 505528 437912
rect 505562 437878 506316 437912
rect 506350 437878 506416 437912
rect 506450 437878 506516 437912
rect 506550 437878 506616 437912
rect 506650 437878 506716 437912
rect 506750 437878 506816 437912
rect 506850 437878 507604 437912
rect 507638 437878 507704 437912
rect 507738 437878 507804 437912
rect 507838 437878 507904 437912
rect 507938 437878 508004 437912
rect 508038 437878 508104 437912
rect 508138 437878 508892 437912
rect 508926 437878 508992 437912
rect 509026 437878 509092 437912
rect 509126 437878 509192 437912
rect 509226 437878 509292 437912
rect 509326 437878 509392 437912
rect 509426 437878 510180 437912
rect 510214 437878 510280 437912
rect 510314 437878 510380 437912
rect 510414 437878 510480 437912
rect 510514 437878 510580 437912
rect 510614 437878 510680 437912
rect 510714 437878 511468 437912
rect 511502 437878 511568 437912
rect 511602 437878 511668 437912
rect 511702 437878 511768 437912
rect 511802 437878 511868 437912
rect 511902 437878 511968 437912
rect 512002 437878 512756 437912
rect 512790 437878 512856 437912
rect 512890 437878 512956 437912
rect 512990 437878 513056 437912
rect 513090 437878 513156 437912
rect 513190 437878 513256 437912
rect 513290 437878 513335 437912
rect 503709 437812 513335 437878
rect 503709 437778 503740 437812
rect 503774 437778 503840 437812
rect 503874 437778 503940 437812
rect 503974 437778 504040 437812
rect 504074 437778 504140 437812
rect 504174 437778 504240 437812
rect 504274 437778 505028 437812
rect 505062 437778 505128 437812
rect 505162 437778 505228 437812
rect 505262 437778 505328 437812
rect 505362 437778 505428 437812
rect 505462 437778 505528 437812
rect 505562 437778 506316 437812
rect 506350 437778 506416 437812
rect 506450 437778 506516 437812
rect 506550 437778 506616 437812
rect 506650 437778 506716 437812
rect 506750 437778 506816 437812
rect 506850 437778 507604 437812
rect 507638 437778 507704 437812
rect 507738 437778 507804 437812
rect 507838 437778 507904 437812
rect 507938 437778 508004 437812
rect 508038 437778 508104 437812
rect 508138 437778 508892 437812
rect 508926 437778 508992 437812
rect 509026 437778 509092 437812
rect 509126 437778 509192 437812
rect 509226 437778 509292 437812
rect 509326 437778 509392 437812
rect 509426 437778 510180 437812
rect 510214 437778 510280 437812
rect 510314 437778 510380 437812
rect 510414 437778 510480 437812
rect 510514 437778 510580 437812
rect 510614 437778 510680 437812
rect 510714 437778 511468 437812
rect 511502 437778 511568 437812
rect 511602 437778 511668 437812
rect 511702 437778 511768 437812
rect 511802 437778 511868 437812
rect 511902 437778 511968 437812
rect 512002 437778 512756 437812
rect 512790 437778 512856 437812
rect 512890 437778 512956 437812
rect 512990 437778 513056 437812
rect 513090 437778 513156 437812
rect 513190 437778 513256 437812
rect 513290 437778 513335 437812
rect 503709 437712 513335 437778
rect 503709 437678 503740 437712
rect 503774 437678 503840 437712
rect 503874 437678 503940 437712
rect 503974 437678 504040 437712
rect 504074 437678 504140 437712
rect 504174 437678 504240 437712
rect 504274 437678 505028 437712
rect 505062 437678 505128 437712
rect 505162 437678 505228 437712
rect 505262 437678 505328 437712
rect 505362 437678 505428 437712
rect 505462 437678 505528 437712
rect 505562 437678 506316 437712
rect 506350 437678 506416 437712
rect 506450 437678 506516 437712
rect 506550 437678 506616 437712
rect 506650 437678 506716 437712
rect 506750 437678 506816 437712
rect 506850 437678 507604 437712
rect 507638 437678 507704 437712
rect 507738 437678 507804 437712
rect 507838 437678 507904 437712
rect 507938 437678 508004 437712
rect 508038 437678 508104 437712
rect 508138 437678 508892 437712
rect 508926 437678 508992 437712
rect 509026 437678 509092 437712
rect 509126 437678 509192 437712
rect 509226 437678 509292 437712
rect 509326 437678 509392 437712
rect 509426 437678 510180 437712
rect 510214 437678 510280 437712
rect 510314 437678 510380 437712
rect 510414 437678 510480 437712
rect 510514 437678 510580 437712
rect 510614 437678 510680 437712
rect 510714 437678 511468 437712
rect 511502 437678 511568 437712
rect 511602 437678 511668 437712
rect 511702 437678 511768 437712
rect 511802 437678 511868 437712
rect 511902 437678 511968 437712
rect 512002 437678 512756 437712
rect 512790 437678 512856 437712
rect 512890 437678 512956 437712
rect 512990 437678 513056 437712
rect 513090 437678 513156 437712
rect 513190 437678 513256 437712
rect 513290 437678 513335 437712
rect 503709 437612 513335 437678
rect 500384 437540 501444 437580
rect 500384 437440 500418 437540
rect 500518 437440 500642 437540
rect 500742 437440 500866 437540
rect 500966 437440 501090 437540
rect 501190 437440 501314 437540
rect 501414 437440 501444 437540
rect 500384 437316 501444 437440
rect 500384 437216 500418 437316
rect 500518 437216 500642 437316
rect 500742 437216 500866 437316
rect 500966 437216 501090 437316
rect 501190 437216 501314 437316
rect 501414 437216 501444 437316
rect 500384 437092 501444 437216
rect 500384 436992 500418 437092
rect 500518 436992 500642 437092
rect 500742 436992 500866 437092
rect 500966 436992 501090 437092
rect 501190 436992 501314 437092
rect 501414 436992 501444 437092
rect 500384 436868 501444 436992
rect 500384 436768 500418 436868
rect 500518 436768 500642 436868
rect 500742 436768 500866 436868
rect 500966 436768 501090 436868
rect 501190 436768 501314 436868
rect 501414 436768 501444 436868
rect 500384 436644 501444 436768
rect 500384 436544 500418 436644
rect 500518 436544 500642 436644
rect 500742 436544 500866 436644
rect 500966 436544 501090 436644
rect 501190 436544 501314 436644
rect 501414 436544 501444 436644
rect 500384 436420 501444 436544
rect 500384 436320 500418 436420
rect 500518 436320 500642 436420
rect 500742 436320 500866 436420
rect 500966 436320 501090 436420
rect 501190 436320 501314 436420
rect 501414 436320 501444 436420
rect 500384 436196 501444 436320
rect 500384 436096 500418 436196
rect 500518 436096 500642 436196
rect 500742 436096 500866 436196
rect 500966 436096 501090 436196
rect 501190 436096 501314 436196
rect 501414 436096 501444 436196
rect 500384 435972 501444 436096
rect 500384 435872 500418 435972
rect 500518 435872 500642 435972
rect 500742 435872 500866 435972
rect 500966 435872 501090 435972
rect 501190 435872 501314 435972
rect 501414 435872 501444 435972
rect 500384 435748 501444 435872
rect 500384 435648 500418 435748
rect 500518 435648 500642 435748
rect 500742 435648 500866 435748
rect 500966 435648 501090 435748
rect 501190 435648 501314 435748
rect 501414 435648 501444 435748
rect 500384 435524 501444 435648
rect 500384 435424 500418 435524
rect 500518 435424 500642 435524
rect 500742 435424 500866 435524
rect 500966 435424 501090 435524
rect 501190 435424 501314 435524
rect 501414 435424 501444 435524
rect 500384 435300 501444 435424
rect 500384 435200 500418 435300
rect 500518 435200 500642 435300
rect 500742 435200 500866 435300
rect 500966 435200 501090 435300
rect 501190 435200 501314 435300
rect 501414 435200 501444 435300
rect 500384 435076 501444 435200
rect 500384 434976 500418 435076
rect 500518 434976 500642 435076
rect 500742 434976 500866 435076
rect 500966 434976 501090 435076
rect 501190 434976 501314 435076
rect 501414 434976 501444 435076
rect 500384 434852 501444 434976
rect 500384 434752 500418 434852
rect 500518 434752 500642 434852
rect 500742 434752 500866 434852
rect 500966 434752 501090 434852
rect 501190 434752 501314 434852
rect 501414 434752 501444 434852
rect 500384 434628 501444 434752
rect 500384 434528 500418 434628
rect 500518 434528 500642 434628
rect 500742 434528 500866 434628
rect 500966 434528 501090 434628
rect 501190 434528 501314 434628
rect 501414 434528 501444 434628
rect 500384 434404 501444 434528
rect 500384 434304 500418 434404
rect 500518 434304 500642 434404
rect 500742 434304 500866 434404
rect 500966 434304 501090 434404
rect 501190 434304 501314 434404
rect 501414 434304 501444 434404
rect 500384 434180 501444 434304
rect 500384 434080 500418 434180
rect 500518 434080 500642 434180
rect 500742 434080 500866 434180
rect 500966 434080 501090 434180
rect 501190 434080 501314 434180
rect 501414 434080 501444 434180
rect 500384 433956 501444 434080
rect 500384 433856 500418 433956
rect 500518 433856 500642 433956
rect 500742 433856 500866 433956
rect 500966 433856 501090 433956
rect 501190 433856 501314 433956
rect 501414 433856 501444 433956
rect 500384 433732 501444 433856
rect 500384 433632 500418 433732
rect 500518 433632 500642 433732
rect 500742 433632 500866 433732
rect 500966 433632 501090 433732
rect 501190 433632 501314 433732
rect 501414 433632 501444 433732
rect 500384 433508 501444 433632
rect 500384 433408 500418 433508
rect 500518 433408 500642 433508
rect 500742 433408 500866 433508
rect 500966 433408 501090 433508
rect 501190 433408 501314 433508
rect 501414 433408 501444 433508
rect 500384 433284 501444 433408
rect 500384 433184 500418 433284
rect 500518 433184 500642 433284
rect 500742 433184 500866 433284
rect 500966 433184 501090 433284
rect 501190 433184 501314 433284
rect 501414 433184 501444 433284
rect 500384 433060 501444 433184
rect 500384 432960 500418 433060
rect 500518 432960 500642 433060
rect 500742 432960 500866 433060
rect 500966 432960 501090 433060
rect 501190 432960 501314 433060
rect 501414 432960 501444 433060
rect 500384 432836 501444 432960
rect 500384 432736 500418 432836
rect 500518 432736 500642 432836
rect 500742 432736 500866 432836
rect 500966 432736 501090 432836
rect 501190 432736 501314 432836
rect 501414 432736 501444 432836
rect 500384 432612 501444 432736
rect 500384 432512 500418 432612
rect 500518 432512 500642 432612
rect 500742 432512 500866 432612
rect 500966 432512 501090 432612
rect 501190 432512 501314 432612
rect 501414 432512 501444 432612
rect 500384 432388 501444 432512
rect 500384 432288 500418 432388
rect 500518 432288 500642 432388
rect 500742 432288 500866 432388
rect 500966 432288 501090 432388
rect 501190 432288 501314 432388
rect 501414 432288 501444 432388
rect 503709 437578 503740 437612
rect 503774 437578 503840 437612
rect 503874 437578 503940 437612
rect 503974 437578 504040 437612
rect 504074 437578 504140 437612
rect 504174 437578 504240 437612
rect 504274 437578 505028 437612
rect 505062 437578 505128 437612
rect 505162 437578 505228 437612
rect 505262 437578 505328 437612
rect 505362 437578 505428 437612
rect 505462 437578 505528 437612
rect 505562 437578 506316 437612
rect 506350 437578 506416 437612
rect 506450 437578 506516 437612
rect 506550 437578 506616 437612
rect 506650 437578 506716 437612
rect 506750 437578 506816 437612
rect 506850 437578 507604 437612
rect 507638 437578 507704 437612
rect 507738 437578 507804 437612
rect 507838 437578 507904 437612
rect 507938 437578 508004 437612
rect 508038 437578 508104 437612
rect 508138 437578 508892 437612
rect 508926 437578 508992 437612
rect 509026 437578 509092 437612
rect 509126 437578 509192 437612
rect 509226 437578 509292 437612
rect 509326 437578 509392 437612
rect 509426 437578 510180 437612
rect 510214 437578 510280 437612
rect 510314 437578 510380 437612
rect 510414 437578 510480 437612
rect 510514 437578 510580 437612
rect 510614 437578 510680 437612
rect 510714 437578 511468 437612
rect 511502 437578 511568 437612
rect 511602 437578 511668 437612
rect 511702 437578 511768 437612
rect 511802 437578 511868 437612
rect 511902 437578 511968 437612
rect 512002 437578 512756 437612
rect 512790 437578 512856 437612
rect 512890 437578 512956 437612
rect 512990 437578 513056 437612
rect 513090 437578 513156 437612
rect 513190 437578 513256 437612
rect 513290 437578 513335 437612
rect 503709 436848 513335 437578
rect 503709 436796 503716 436848
rect 503768 436824 503820 436848
rect 503872 436824 503924 436848
rect 503774 436796 503820 436824
rect 503874 436796 503924 436824
rect 503976 436796 504028 436848
rect 504080 436796 504132 436848
rect 504184 436796 504236 436848
rect 504288 436824 513335 436848
rect 504288 436796 505028 436824
rect 503709 436790 503740 436796
rect 503774 436790 503840 436796
rect 503874 436790 503940 436796
rect 503974 436790 504040 436796
rect 504074 436790 504140 436796
rect 504174 436790 504240 436796
rect 504274 436790 505028 436796
rect 505062 436790 505128 436824
rect 505162 436790 505228 436824
rect 505262 436790 505328 436824
rect 505362 436790 505428 436824
rect 505462 436790 505528 436824
rect 505562 436790 506316 436824
rect 506350 436790 506416 436824
rect 506450 436790 506516 436824
rect 506550 436790 506616 436824
rect 506650 436790 506716 436824
rect 506750 436790 506816 436824
rect 506850 436790 507604 436824
rect 507638 436790 507704 436824
rect 507738 436790 507804 436824
rect 507838 436790 507904 436824
rect 507938 436790 508004 436824
rect 508038 436790 508104 436824
rect 508138 436790 508892 436824
rect 508926 436790 508992 436824
rect 509026 436790 509092 436824
rect 509126 436790 509192 436824
rect 509226 436790 509292 436824
rect 509326 436790 509392 436824
rect 509426 436790 510180 436824
rect 510214 436790 510280 436824
rect 510314 436790 510380 436824
rect 510414 436790 510480 436824
rect 510514 436790 510580 436824
rect 510614 436790 510680 436824
rect 510714 436790 511468 436824
rect 511502 436790 511568 436824
rect 511602 436790 511668 436824
rect 511702 436790 511768 436824
rect 511802 436790 511868 436824
rect 511902 436790 511968 436824
rect 512002 436790 512756 436824
rect 512790 436790 512856 436824
rect 512890 436790 512956 436824
rect 512990 436790 513056 436824
rect 513090 436790 513156 436824
rect 513190 436790 513256 436824
rect 513290 436790 513335 436824
rect 503709 436744 513335 436790
rect 503709 436692 503716 436744
rect 503768 436724 503820 436744
rect 503872 436724 503924 436744
rect 503774 436692 503820 436724
rect 503874 436692 503924 436724
rect 503976 436692 504028 436744
rect 504080 436692 504132 436744
rect 504184 436692 504236 436744
rect 504288 436724 513335 436744
rect 504288 436692 505028 436724
rect 503709 436690 503740 436692
rect 503774 436690 503840 436692
rect 503874 436690 503940 436692
rect 503974 436690 504040 436692
rect 504074 436690 504140 436692
rect 504174 436690 504240 436692
rect 504274 436690 505028 436692
rect 505062 436690 505128 436724
rect 505162 436690 505228 436724
rect 505262 436690 505328 436724
rect 505362 436690 505428 436724
rect 505462 436690 505528 436724
rect 505562 436690 506316 436724
rect 506350 436690 506416 436724
rect 506450 436690 506516 436724
rect 506550 436690 506616 436724
rect 506650 436690 506716 436724
rect 506750 436690 506816 436724
rect 506850 436690 507604 436724
rect 507638 436690 507704 436724
rect 507738 436690 507804 436724
rect 507838 436690 507904 436724
rect 507938 436690 508004 436724
rect 508038 436690 508104 436724
rect 508138 436690 508892 436724
rect 508926 436690 508992 436724
rect 509026 436690 509092 436724
rect 509126 436690 509192 436724
rect 509226 436690 509292 436724
rect 509326 436690 509392 436724
rect 509426 436690 510180 436724
rect 510214 436690 510280 436724
rect 510314 436690 510380 436724
rect 510414 436690 510480 436724
rect 510514 436690 510580 436724
rect 510614 436690 510680 436724
rect 510714 436690 511468 436724
rect 511502 436690 511568 436724
rect 511602 436690 511668 436724
rect 511702 436690 511768 436724
rect 511802 436690 511868 436724
rect 511902 436690 511968 436724
rect 512002 436690 512756 436724
rect 512790 436690 512856 436724
rect 512890 436690 512956 436724
rect 512990 436690 513056 436724
rect 513090 436690 513156 436724
rect 513190 436690 513256 436724
rect 513290 436690 513335 436724
rect 503709 436640 513335 436690
rect 503709 436588 503716 436640
rect 503768 436624 503820 436640
rect 503872 436624 503924 436640
rect 503774 436590 503820 436624
rect 503874 436590 503924 436624
rect 503768 436588 503820 436590
rect 503872 436588 503924 436590
rect 503976 436588 504028 436640
rect 504080 436588 504132 436640
rect 504184 436588 504236 436640
rect 504288 436624 513335 436640
rect 504288 436590 505028 436624
rect 505062 436590 505128 436624
rect 505162 436590 505228 436624
rect 505262 436590 505328 436624
rect 505362 436590 505428 436624
rect 505462 436590 505528 436624
rect 505562 436590 506316 436624
rect 506350 436590 506416 436624
rect 506450 436590 506516 436624
rect 506550 436590 506616 436624
rect 506650 436590 506716 436624
rect 506750 436590 506816 436624
rect 506850 436590 507604 436624
rect 507638 436590 507704 436624
rect 507738 436590 507804 436624
rect 507838 436590 507904 436624
rect 507938 436590 508004 436624
rect 508038 436590 508104 436624
rect 508138 436590 508892 436624
rect 508926 436590 508992 436624
rect 509026 436590 509092 436624
rect 509126 436590 509192 436624
rect 509226 436590 509292 436624
rect 509326 436590 509392 436624
rect 509426 436590 510180 436624
rect 510214 436590 510280 436624
rect 510314 436590 510380 436624
rect 510414 436590 510480 436624
rect 510514 436590 510580 436624
rect 510614 436590 510680 436624
rect 510714 436590 511468 436624
rect 511502 436590 511568 436624
rect 511602 436590 511668 436624
rect 511702 436590 511768 436624
rect 511802 436590 511868 436624
rect 511902 436590 511968 436624
rect 512002 436590 512756 436624
rect 512790 436590 512856 436624
rect 512890 436590 512956 436624
rect 512990 436590 513056 436624
rect 513090 436590 513156 436624
rect 513190 436590 513256 436624
rect 513290 436590 513335 436624
rect 504288 436588 513335 436590
rect 503709 436536 513335 436588
rect 503709 436484 503716 436536
rect 503768 436524 503820 436536
rect 503872 436524 503924 436536
rect 503774 436490 503820 436524
rect 503874 436490 503924 436524
rect 503768 436484 503820 436490
rect 503872 436484 503924 436490
rect 503976 436484 504028 436536
rect 504080 436484 504132 436536
rect 504184 436484 504236 436536
rect 504288 436524 513335 436536
rect 504288 436490 505028 436524
rect 505062 436490 505128 436524
rect 505162 436490 505228 436524
rect 505262 436490 505328 436524
rect 505362 436490 505428 436524
rect 505462 436490 505528 436524
rect 505562 436490 506316 436524
rect 506350 436490 506416 436524
rect 506450 436490 506516 436524
rect 506550 436490 506616 436524
rect 506650 436490 506716 436524
rect 506750 436490 506816 436524
rect 506850 436490 507604 436524
rect 507638 436490 507704 436524
rect 507738 436490 507804 436524
rect 507838 436490 507904 436524
rect 507938 436490 508004 436524
rect 508038 436490 508104 436524
rect 508138 436490 508892 436524
rect 508926 436490 508992 436524
rect 509026 436490 509092 436524
rect 509126 436490 509192 436524
rect 509226 436490 509292 436524
rect 509326 436490 509392 436524
rect 509426 436490 510180 436524
rect 510214 436490 510280 436524
rect 510314 436490 510380 436524
rect 510414 436490 510480 436524
rect 510514 436490 510580 436524
rect 510614 436490 510680 436524
rect 510714 436490 511468 436524
rect 511502 436490 511568 436524
rect 511602 436490 511668 436524
rect 511702 436490 511768 436524
rect 511802 436490 511868 436524
rect 511902 436490 511968 436524
rect 512002 436490 512756 436524
rect 512790 436490 512856 436524
rect 512890 436490 512956 436524
rect 512990 436490 513056 436524
rect 513090 436490 513156 436524
rect 513190 436490 513256 436524
rect 513290 436490 513335 436524
rect 504288 436484 513335 436490
rect 503709 436432 513335 436484
rect 503709 436380 503716 436432
rect 503768 436424 503820 436432
rect 503872 436424 503924 436432
rect 503774 436390 503820 436424
rect 503874 436390 503924 436424
rect 503768 436380 503820 436390
rect 503872 436380 503924 436390
rect 503976 436380 504028 436432
rect 504080 436380 504132 436432
rect 504184 436380 504236 436432
rect 504288 436424 513335 436432
rect 504288 436390 505028 436424
rect 505062 436390 505128 436424
rect 505162 436390 505228 436424
rect 505262 436390 505328 436424
rect 505362 436390 505428 436424
rect 505462 436390 505528 436424
rect 505562 436390 506316 436424
rect 506350 436390 506416 436424
rect 506450 436390 506516 436424
rect 506550 436390 506616 436424
rect 506650 436390 506716 436424
rect 506750 436390 506816 436424
rect 506850 436390 507604 436424
rect 507638 436390 507704 436424
rect 507738 436390 507804 436424
rect 507838 436390 507904 436424
rect 507938 436390 508004 436424
rect 508038 436390 508104 436424
rect 508138 436390 508892 436424
rect 508926 436390 508992 436424
rect 509026 436390 509092 436424
rect 509126 436390 509192 436424
rect 509226 436390 509292 436424
rect 509326 436390 509392 436424
rect 509426 436390 510180 436424
rect 510214 436390 510280 436424
rect 510314 436390 510380 436424
rect 510414 436390 510480 436424
rect 510514 436390 510580 436424
rect 510614 436390 510680 436424
rect 510714 436390 511468 436424
rect 511502 436390 511568 436424
rect 511602 436390 511668 436424
rect 511702 436390 511768 436424
rect 511802 436390 511868 436424
rect 511902 436390 511968 436424
rect 512002 436390 512756 436424
rect 512790 436390 512856 436424
rect 512890 436390 512956 436424
rect 512990 436390 513056 436424
rect 513090 436390 513156 436424
rect 513190 436390 513256 436424
rect 513290 436390 513335 436424
rect 504288 436380 513335 436390
rect 503709 436328 513335 436380
rect 503709 436276 503716 436328
rect 503768 436324 503820 436328
rect 503872 436324 503924 436328
rect 503774 436290 503820 436324
rect 503874 436290 503924 436324
rect 503768 436276 503820 436290
rect 503872 436276 503924 436290
rect 503976 436276 504028 436328
rect 504080 436276 504132 436328
rect 504184 436276 504236 436328
rect 504288 436324 513335 436328
rect 504288 436290 505028 436324
rect 505062 436290 505128 436324
rect 505162 436290 505228 436324
rect 505262 436290 505328 436324
rect 505362 436290 505428 436324
rect 505462 436290 505528 436324
rect 505562 436290 506316 436324
rect 506350 436290 506416 436324
rect 506450 436290 506516 436324
rect 506550 436290 506616 436324
rect 506650 436290 506716 436324
rect 506750 436290 506816 436324
rect 506850 436290 507604 436324
rect 507638 436290 507704 436324
rect 507738 436290 507804 436324
rect 507838 436290 507904 436324
rect 507938 436290 508004 436324
rect 508038 436290 508104 436324
rect 508138 436290 508892 436324
rect 508926 436290 508992 436324
rect 509026 436290 509092 436324
rect 509126 436290 509192 436324
rect 509226 436290 509292 436324
rect 509326 436290 509392 436324
rect 509426 436290 510180 436324
rect 510214 436290 510280 436324
rect 510314 436290 510380 436324
rect 510414 436290 510480 436324
rect 510514 436290 510580 436324
rect 510614 436290 510680 436324
rect 510714 436290 511468 436324
rect 511502 436290 511568 436324
rect 511602 436290 511668 436324
rect 511702 436290 511768 436324
rect 511802 436290 511868 436324
rect 511902 436290 511968 436324
rect 512002 436290 512756 436324
rect 512790 436290 512856 436324
rect 512890 436290 512956 436324
rect 512990 436290 513056 436324
rect 513090 436290 513156 436324
rect 513190 436290 513256 436324
rect 513290 436290 513335 436324
rect 504288 436276 513335 436290
rect 503709 436245 513335 436276
rect 503709 435536 508183 436245
rect 503709 435502 503740 435536
rect 503774 435502 503840 435536
rect 503874 435502 503940 435536
rect 503974 435502 504040 435536
rect 504074 435502 504140 435536
rect 504174 435502 504240 435536
rect 504274 435502 505028 435536
rect 505062 435502 505128 435536
rect 505162 435502 505228 435536
rect 505262 435502 505328 435536
rect 505362 435502 505428 435536
rect 505462 435502 505528 435536
rect 505562 435502 506316 435536
rect 506350 435502 506416 435536
rect 506450 435502 506516 435536
rect 506550 435502 506616 435536
rect 506650 435502 506716 435536
rect 506750 435502 506816 435536
rect 506850 435502 507604 435536
rect 507638 435502 507704 435536
rect 507738 435502 507804 435536
rect 507838 435502 507904 435536
rect 507938 435502 508004 435536
rect 508038 435502 508104 435536
rect 508138 435502 508183 435536
rect 503709 435436 508183 435502
rect 503709 435402 503740 435436
rect 503774 435402 503840 435436
rect 503874 435402 503940 435436
rect 503974 435402 504040 435436
rect 504074 435402 504140 435436
rect 504174 435402 504240 435436
rect 504274 435402 505028 435436
rect 505062 435402 505128 435436
rect 505162 435402 505228 435436
rect 505262 435402 505328 435436
rect 505362 435402 505428 435436
rect 505462 435402 505528 435436
rect 505562 435402 506316 435436
rect 506350 435402 506416 435436
rect 506450 435402 506516 435436
rect 506550 435402 506616 435436
rect 506650 435402 506716 435436
rect 506750 435402 506816 435436
rect 506850 435402 507604 435436
rect 507638 435402 507704 435436
rect 507738 435402 507804 435436
rect 507838 435402 507904 435436
rect 507938 435402 508004 435436
rect 508038 435402 508104 435436
rect 508138 435402 508183 435436
rect 503709 435336 508183 435402
rect 503709 435302 503740 435336
rect 503774 435302 503840 435336
rect 503874 435302 503940 435336
rect 503974 435302 504040 435336
rect 504074 435302 504140 435336
rect 504174 435302 504240 435336
rect 504274 435302 505028 435336
rect 505062 435302 505128 435336
rect 505162 435302 505228 435336
rect 505262 435302 505328 435336
rect 505362 435302 505428 435336
rect 505462 435302 505528 435336
rect 505562 435302 506316 435336
rect 506350 435302 506416 435336
rect 506450 435302 506516 435336
rect 506550 435302 506616 435336
rect 506650 435302 506716 435336
rect 506750 435302 506816 435336
rect 506850 435302 507604 435336
rect 507638 435302 507704 435336
rect 507738 435302 507804 435336
rect 507838 435302 507904 435336
rect 507938 435302 508004 435336
rect 508038 435302 508104 435336
rect 508138 435302 508183 435336
rect 503709 435236 508183 435302
rect 503709 435202 503740 435236
rect 503774 435202 503840 435236
rect 503874 435202 503940 435236
rect 503974 435202 504040 435236
rect 504074 435202 504140 435236
rect 504174 435202 504240 435236
rect 504274 435202 505028 435236
rect 505062 435202 505128 435236
rect 505162 435202 505228 435236
rect 505262 435202 505328 435236
rect 505362 435202 505428 435236
rect 505462 435202 505528 435236
rect 505562 435202 506316 435236
rect 506350 435202 506416 435236
rect 506450 435202 506516 435236
rect 506550 435202 506616 435236
rect 506650 435202 506716 435236
rect 506750 435202 506816 435236
rect 506850 435202 507604 435236
rect 507638 435202 507704 435236
rect 507738 435202 507804 435236
rect 507838 435202 507904 435236
rect 507938 435202 508004 435236
rect 508038 435202 508104 435236
rect 508138 435202 508183 435236
rect 503709 435136 508183 435202
rect 503709 435102 503740 435136
rect 503774 435102 503840 435136
rect 503874 435102 503940 435136
rect 503974 435102 504040 435136
rect 504074 435102 504140 435136
rect 504174 435102 504240 435136
rect 504274 435102 505028 435136
rect 505062 435102 505128 435136
rect 505162 435102 505228 435136
rect 505262 435102 505328 435136
rect 505362 435102 505428 435136
rect 505462 435102 505528 435136
rect 505562 435102 506316 435136
rect 506350 435102 506416 435136
rect 506450 435102 506516 435136
rect 506550 435102 506616 435136
rect 506650 435102 506716 435136
rect 506750 435102 506816 435136
rect 506850 435102 507604 435136
rect 507638 435102 507704 435136
rect 507738 435102 507804 435136
rect 507838 435102 507904 435136
rect 507938 435102 508004 435136
rect 508038 435102 508104 435136
rect 508138 435102 508183 435136
rect 503709 435036 508183 435102
rect 503709 435002 503740 435036
rect 503774 435002 503840 435036
rect 503874 435002 503940 435036
rect 503974 435002 504040 435036
rect 504074 435002 504140 435036
rect 504174 435002 504240 435036
rect 504274 435002 505028 435036
rect 505062 435002 505128 435036
rect 505162 435002 505228 435036
rect 505262 435002 505328 435036
rect 505362 435002 505428 435036
rect 505462 435002 505528 435036
rect 505562 435002 506316 435036
rect 506350 435002 506416 435036
rect 506450 435002 506516 435036
rect 506550 435002 506616 435036
rect 506650 435002 506716 435036
rect 506750 435002 506816 435036
rect 506850 435002 507604 435036
rect 507638 435002 507704 435036
rect 507738 435002 507804 435036
rect 507838 435002 507904 435036
rect 507938 435002 508004 435036
rect 508038 435002 508104 435036
rect 508138 435002 508183 435036
rect 503709 434279 508183 435002
rect 508861 435560 509471 435567
rect 508861 435508 508868 435560
rect 508920 435536 508972 435560
rect 509024 435536 509076 435560
rect 508926 435508 508972 435536
rect 509026 435508 509076 435536
rect 509128 435508 509180 435560
rect 509232 435508 509284 435560
rect 509336 435508 509388 435560
rect 509440 435508 509471 435560
rect 508861 435502 508892 435508
rect 508926 435502 508992 435508
rect 509026 435502 509092 435508
rect 509126 435502 509192 435508
rect 509226 435502 509292 435508
rect 509326 435502 509392 435508
rect 509426 435502 509471 435508
rect 508861 435456 509471 435502
rect 508861 435404 508868 435456
rect 508920 435436 508972 435456
rect 509024 435436 509076 435456
rect 508926 435404 508972 435436
rect 509026 435404 509076 435436
rect 509128 435404 509180 435456
rect 509232 435404 509284 435456
rect 509336 435404 509388 435456
rect 509440 435404 509471 435456
rect 508861 435402 508892 435404
rect 508926 435402 508992 435404
rect 509026 435402 509092 435404
rect 509126 435402 509192 435404
rect 509226 435402 509292 435404
rect 509326 435402 509392 435404
rect 509426 435402 509471 435404
rect 508861 435352 509471 435402
rect 508861 435300 508868 435352
rect 508920 435336 508972 435352
rect 509024 435336 509076 435352
rect 508926 435302 508972 435336
rect 509026 435302 509076 435336
rect 508920 435300 508972 435302
rect 509024 435300 509076 435302
rect 509128 435300 509180 435352
rect 509232 435300 509284 435352
rect 509336 435300 509388 435352
rect 509440 435300 509471 435352
rect 508861 435248 509471 435300
rect 508861 435196 508868 435248
rect 508920 435236 508972 435248
rect 509024 435236 509076 435248
rect 508926 435202 508972 435236
rect 509026 435202 509076 435236
rect 508920 435196 508972 435202
rect 509024 435196 509076 435202
rect 509128 435196 509180 435248
rect 509232 435196 509284 435248
rect 509336 435196 509388 435248
rect 509440 435196 509471 435248
rect 508861 435144 509471 435196
rect 508861 435092 508868 435144
rect 508920 435136 508972 435144
rect 509024 435136 509076 435144
rect 508926 435102 508972 435136
rect 509026 435102 509076 435136
rect 508920 435092 508972 435102
rect 509024 435092 509076 435102
rect 509128 435092 509180 435144
rect 509232 435092 509284 435144
rect 509336 435092 509388 435144
rect 509440 435092 509471 435144
rect 508861 435040 509471 435092
rect 508861 434988 508868 435040
rect 508920 435036 508972 435040
rect 509024 435036 509076 435040
rect 508926 435002 508972 435036
rect 509026 435002 509076 435036
rect 508920 434988 508972 435002
rect 509024 434988 509076 435002
rect 509128 434988 509180 435040
rect 509232 434988 509284 435040
rect 509336 434988 509388 435040
rect 509440 434988 509471 435040
rect 508861 434957 509471 434988
rect 510149 435536 513335 436245
rect 510149 435502 510180 435536
rect 510214 435502 510280 435536
rect 510314 435502 510380 435536
rect 510414 435502 510480 435536
rect 510514 435502 510580 435536
rect 510614 435502 510680 435536
rect 510714 435502 511468 435536
rect 511502 435502 511568 435536
rect 511602 435502 511668 435536
rect 511702 435502 511768 435536
rect 511802 435502 511868 435536
rect 511902 435502 511968 435536
rect 512002 435502 512756 435536
rect 512790 435502 512856 435536
rect 512890 435502 512956 435536
rect 512990 435502 513056 435536
rect 513090 435502 513156 435536
rect 513190 435502 513256 435536
rect 513290 435502 513335 435536
rect 510149 435436 513335 435502
rect 510149 435402 510180 435436
rect 510214 435402 510280 435436
rect 510314 435402 510380 435436
rect 510414 435402 510480 435436
rect 510514 435402 510580 435436
rect 510614 435402 510680 435436
rect 510714 435402 511468 435436
rect 511502 435402 511568 435436
rect 511602 435402 511668 435436
rect 511702 435402 511768 435436
rect 511802 435402 511868 435436
rect 511902 435402 511968 435436
rect 512002 435402 512756 435436
rect 512790 435402 512856 435436
rect 512890 435402 512956 435436
rect 512990 435402 513056 435436
rect 513090 435402 513156 435436
rect 513190 435402 513256 435436
rect 513290 435402 513335 435436
rect 510149 435336 513335 435402
rect 510149 435302 510180 435336
rect 510214 435302 510280 435336
rect 510314 435302 510380 435336
rect 510414 435302 510480 435336
rect 510514 435302 510580 435336
rect 510614 435302 510680 435336
rect 510714 435302 511468 435336
rect 511502 435302 511568 435336
rect 511602 435302 511668 435336
rect 511702 435302 511768 435336
rect 511802 435302 511868 435336
rect 511902 435302 511968 435336
rect 512002 435302 512756 435336
rect 512790 435302 512856 435336
rect 512890 435302 512956 435336
rect 512990 435302 513056 435336
rect 513090 435302 513156 435336
rect 513190 435302 513256 435336
rect 513290 435302 513335 435336
rect 510149 435236 513335 435302
rect 510149 435202 510180 435236
rect 510214 435202 510280 435236
rect 510314 435202 510380 435236
rect 510414 435202 510480 435236
rect 510514 435202 510580 435236
rect 510614 435202 510680 435236
rect 510714 435202 511468 435236
rect 511502 435202 511568 435236
rect 511602 435202 511668 435236
rect 511702 435202 511768 435236
rect 511802 435202 511868 435236
rect 511902 435202 511968 435236
rect 512002 435202 512756 435236
rect 512790 435202 512856 435236
rect 512890 435202 512956 435236
rect 512990 435202 513056 435236
rect 513090 435202 513156 435236
rect 513190 435202 513256 435236
rect 513290 435202 513335 435236
rect 510149 435136 513335 435202
rect 510149 435102 510180 435136
rect 510214 435102 510280 435136
rect 510314 435102 510380 435136
rect 510414 435102 510480 435136
rect 510514 435102 510580 435136
rect 510614 435102 510680 435136
rect 510714 435102 511468 435136
rect 511502 435102 511568 435136
rect 511602 435102 511668 435136
rect 511702 435102 511768 435136
rect 511802 435102 511868 435136
rect 511902 435102 511968 435136
rect 512002 435102 512756 435136
rect 512790 435102 512856 435136
rect 512890 435102 512956 435136
rect 512990 435102 513056 435136
rect 513090 435102 513156 435136
rect 513190 435102 513256 435136
rect 513290 435102 513335 435136
rect 510149 435036 513335 435102
rect 510149 435002 510180 435036
rect 510214 435002 510280 435036
rect 510314 435002 510380 435036
rect 510414 435002 510480 435036
rect 510514 435002 510580 435036
rect 510614 435002 510680 435036
rect 510714 435002 511468 435036
rect 511502 435002 511568 435036
rect 511602 435002 511668 435036
rect 511702 435002 511768 435036
rect 511802 435002 511868 435036
rect 511902 435002 511968 435036
rect 512002 435002 512756 435036
rect 512790 435002 512856 435036
rect 512890 435002 512956 435036
rect 512990 435002 513056 435036
rect 513090 435002 513156 435036
rect 513190 435002 513256 435036
rect 513290 435002 513335 435036
rect 510149 434279 513335 435002
rect 503709 434248 513335 434279
rect 503709 434214 503740 434248
rect 503774 434214 503840 434248
rect 503874 434214 503940 434248
rect 503974 434214 504040 434248
rect 504074 434214 504140 434248
rect 504174 434214 504240 434248
rect 504274 434214 505028 434248
rect 505062 434214 505128 434248
rect 505162 434214 505228 434248
rect 505262 434214 505328 434248
rect 505362 434214 505428 434248
rect 505462 434214 505528 434248
rect 505562 434214 506316 434248
rect 506350 434214 506416 434248
rect 506450 434214 506516 434248
rect 506550 434214 506616 434248
rect 506650 434214 506716 434248
rect 506750 434214 506816 434248
rect 506850 434214 507604 434248
rect 507638 434214 507704 434248
rect 507738 434214 507804 434248
rect 507838 434214 507904 434248
rect 507938 434214 508004 434248
rect 508038 434214 508104 434248
rect 508138 434214 508892 434248
rect 508926 434214 508992 434248
rect 509026 434214 509092 434248
rect 509126 434214 509192 434248
rect 509226 434214 509292 434248
rect 509326 434214 509392 434248
rect 509426 434214 510180 434248
rect 510214 434214 510280 434248
rect 510314 434214 510380 434248
rect 510414 434214 510480 434248
rect 510514 434214 510580 434248
rect 510614 434214 510680 434248
rect 510714 434214 511468 434248
rect 511502 434214 511568 434248
rect 511602 434214 511668 434248
rect 511702 434214 511768 434248
rect 511802 434214 511868 434248
rect 511902 434214 511968 434248
rect 512002 434214 512756 434248
rect 512790 434214 512856 434248
rect 512890 434214 512956 434248
rect 512990 434214 513056 434248
rect 513090 434214 513156 434248
rect 513190 434214 513256 434248
rect 513290 434214 513335 434248
rect 503709 434148 513335 434214
rect 503709 434114 503740 434148
rect 503774 434114 503840 434148
rect 503874 434114 503940 434148
rect 503974 434114 504040 434148
rect 504074 434114 504140 434148
rect 504174 434114 504240 434148
rect 504274 434114 505028 434148
rect 505062 434114 505128 434148
rect 505162 434114 505228 434148
rect 505262 434114 505328 434148
rect 505362 434114 505428 434148
rect 505462 434114 505528 434148
rect 505562 434114 506316 434148
rect 506350 434114 506416 434148
rect 506450 434114 506516 434148
rect 506550 434114 506616 434148
rect 506650 434114 506716 434148
rect 506750 434114 506816 434148
rect 506850 434114 507604 434148
rect 507638 434114 507704 434148
rect 507738 434114 507804 434148
rect 507838 434114 507904 434148
rect 507938 434114 508004 434148
rect 508038 434114 508104 434148
rect 508138 434114 508892 434148
rect 508926 434114 508992 434148
rect 509026 434114 509092 434148
rect 509126 434114 509192 434148
rect 509226 434114 509292 434148
rect 509326 434114 509392 434148
rect 509426 434114 510180 434148
rect 510214 434114 510280 434148
rect 510314 434114 510380 434148
rect 510414 434114 510480 434148
rect 510514 434114 510580 434148
rect 510614 434114 510680 434148
rect 510714 434114 511468 434148
rect 511502 434114 511568 434148
rect 511602 434114 511668 434148
rect 511702 434114 511768 434148
rect 511802 434114 511868 434148
rect 511902 434114 511968 434148
rect 512002 434114 512756 434148
rect 512790 434114 512856 434148
rect 512890 434114 512956 434148
rect 512990 434114 513056 434148
rect 513090 434114 513156 434148
rect 513190 434114 513256 434148
rect 513290 434114 513335 434148
rect 503709 434048 513335 434114
rect 503709 434014 503740 434048
rect 503774 434014 503840 434048
rect 503874 434014 503940 434048
rect 503974 434014 504040 434048
rect 504074 434014 504140 434048
rect 504174 434014 504240 434048
rect 504274 434014 505028 434048
rect 505062 434014 505128 434048
rect 505162 434014 505228 434048
rect 505262 434014 505328 434048
rect 505362 434014 505428 434048
rect 505462 434014 505528 434048
rect 505562 434014 506316 434048
rect 506350 434014 506416 434048
rect 506450 434014 506516 434048
rect 506550 434014 506616 434048
rect 506650 434014 506716 434048
rect 506750 434014 506816 434048
rect 506850 434014 507604 434048
rect 507638 434014 507704 434048
rect 507738 434014 507804 434048
rect 507838 434014 507904 434048
rect 507938 434014 508004 434048
rect 508038 434014 508104 434048
rect 508138 434014 508892 434048
rect 508926 434014 508992 434048
rect 509026 434014 509092 434048
rect 509126 434014 509192 434048
rect 509226 434014 509292 434048
rect 509326 434014 509392 434048
rect 509426 434014 510180 434048
rect 510214 434014 510280 434048
rect 510314 434014 510380 434048
rect 510414 434014 510480 434048
rect 510514 434014 510580 434048
rect 510614 434014 510680 434048
rect 510714 434014 511468 434048
rect 511502 434014 511568 434048
rect 511602 434014 511668 434048
rect 511702 434014 511768 434048
rect 511802 434014 511868 434048
rect 511902 434014 511968 434048
rect 512002 434014 512756 434048
rect 512790 434014 512856 434048
rect 512890 434014 512956 434048
rect 512990 434014 513056 434048
rect 513090 434014 513156 434048
rect 513190 434014 513256 434048
rect 513290 434014 513335 434048
rect 503709 433948 513335 434014
rect 503709 433914 503740 433948
rect 503774 433914 503840 433948
rect 503874 433914 503940 433948
rect 503974 433914 504040 433948
rect 504074 433914 504140 433948
rect 504174 433914 504240 433948
rect 504274 433914 505028 433948
rect 505062 433914 505128 433948
rect 505162 433914 505228 433948
rect 505262 433914 505328 433948
rect 505362 433914 505428 433948
rect 505462 433914 505528 433948
rect 505562 433914 506316 433948
rect 506350 433914 506416 433948
rect 506450 433914 506516 433948
rect 506550 433914 506616 433948
rect 506650 433914 506716 433948
rect 506750 433914 506816 433948
rect 506850 433914 507604 433948
rect 507638 433914 507704 433948
rect 507738 433914 507804 433948
rect 507838 433914 507904 433948
rect 507938 433914 508004 433948
rect 508038 433914 508104 433948
rect 508138 433914 508892 433948
rect 508926 433914 508992 433948
rect 509026 433914 509092 433948
rect 509126 433914 509192 433948
rect 509226 433914 509292 433948
rect 509326 433914 509392 433948
rect 509426 433914 510180 433948
rect 510214 433914 510280 433948
rect 510314 433914 510380 433948
rect 510414 433914 510480 433948
rect 510514 433914 510580 433948
rect 510614 433914 510680 433948
rect 510714 433914 511468 433948
rect 511502 433914 511568 433948
rect 511602 433914 511668 433948
rect 511702 433914 511768 433948
rect 511802 433914 511868 433948
rect 511902 433914 511968 433948
rect 512002 433914 512756 433948
rect 512790 433914 512856 433948
rect 512890 433914 512956 433948
rect 512990 433914 513056 433948
rect 513090 433914 513156 433948
rect 513190 433914 513256 433948
rect 513290 433914 513335 433948
rect 503709 433848 513335 433914
rect 503709 433814 503740 433848
rect 503774 433814 503840 433848
rect 503874 433814 503940 433848
rect 503974 433814 504040 433848
rect 504074 433814 504140 433848
rect 504174 433814 504240 433848
rect 504274 433814 505028 433848
rect 505062 433814 505128 433848
rect 505162 433814 505228 433848
rect 505262 433814 505328 433848
rect 505362 433814 505428 433848
rect 505462 433814 505528 433848
rect 505562 433814 506316 433848
rect 506350 433814 506416 433848
rect 506450 433814 506516 433848
rect 506550 433814 506616 433848
rect 506650 433814 506716 433848
rect 506750 433814 506816 433848
rect 506850 433814 507604 433848
rect 507638 433814 507704 433848
rect 507738 433814 507804 433848
rect 507838 433814 507904 433848
rect 507938 433814 508004 433848
rect 508038 433814 508104 433848
rect 508138 433814 508892 433848
rect 508926 433814 508992 433848
rect 509026 433814 509092 433848
rect 509126 433814 509192 433848
rect 509226 433814 509292 433848
rect 509326 433814 509392 433848
rect 509426 433814 510180 433848
rect 510214 433814 510280 433848
rect 510314 433814 510380 433848
rect 510414 433814 510480 433848
rect 510514 433814 510580 433848
rect 510614 433814 510680 433848
rect 510714 433814 511468 433848
rect 511502 433814 511568 433848
rect 511602 433814 511668 433848
rect 511702 433814 511768 433848
rect 511802 433814 511868 433848
rect 511902 433814 511968 433848
rect 512002 433814 512756 433848
rect 512790 433814 512856 433848
rect 512890 433814 512956 433848
rect 512990 433814 513056 433848
rect 513090 433814 513156 433848
rect 513190 433814 513256 433848
rect 513290 433814 513335 433848
rect 503709 433748 513335 433814
rect 503709 433714 503740 433748
rect 503774 433714 503840 433748
rect 503874 433714 503940 433748
rect 503974 433714 504040 433748
rect 504074 433714 504140 433748
rect 504174 433714 504240 433748
rect 504274 433714 505028 433748
rect 505062 433714 505128 433748
rect 505162 433714 505228 433748
rect 505262 433714 505328 433748
rect 505362 433714 505428 433748
rect 505462 433714 505528 433748
rect 505562 433714 506316 433748
rect 506350 433714 506416 433748
rect 506450 433714 506516 433748
rect 506550 433714 506616 433748
rect 506650 433714 506716 433748
rect 506750 433714 506816 433748
rect 506850 433714 507604 433748
rect 507638 433714 507704 433748
rect 507738 433714 507804 433748
rect 507838 433714 507904 433748
rect 507938 433714 508004 433748
rect 508038 433714 508104 433748
rect 508138 433714 508892 433748
rect 508926 433714 508992 433748
rect 509026 433714 509092 433748
rect 509126 433714 509192 433748
rect 509226 433714 509292 433748
rect 509326 433714 509392 433748
rect 509426 433714 510180 433748
rect 510214 433714 510280 433748
rect 510314 433714 510380 433748
rect 510414 433714 510480 433748
rect 510514 433714 510580 433748
rect 510614 433714 510680 433748
rect 510714 433714 511468 433748
rect 511502 433714 511568 433748
rect 511602 433714 511668 433748
rect 511702 433714 511768 433748
rect 511802 433714 511868 433748
rect 511902 433714 511968 433748
rect 512002 433714 512756 433748
rect 512790 433714 512856 433748
rect 512890 433714 512956 433748
rect 512990 433714 513056 433748
rect 513090 433714 513156 433748
rect 513190 433714 513256 433748
rect 513290 433714 513335 433748
rect 503709 432960 513335 433714
rect 503709 432926 503740 432960
rect 503774 432926 503840 432960
rect 503874 432926 503940 432960
rect 503974 432926 504040 432960
rect 504074 432926 504140 432960
rect 504174 432926 504240 432960
rect 504274 432926 505028 432960
rect 505062 432926 505128 432960
rect 505162 432926 505228 432960
rect 505262 432926 505328 432960
rect 505362 432926 505428 432960
rect 505462 432926 505528 432960
rect 505562 432926 506316 432960
rect 506350 432926 506416 432960
rect 506450 432926 506516 432960
rect 506550 432926 506616 432960
rect 506650 432926 506716 432960
rect 506750 432926 506816 432960
rect 506850 432926 507604 432960
rect 507638 432926 507704 432960
rect 507738 432926 507804 432960
rect 507838 432926 507904 432960
rect 507938 432926 508004 432960
rect 508038 432926 508104 432960
rect 508138 432926 508892 432960
rect 508926 432926 508992 432960
rect 509026 432926 509092 432960
rect 509126 432926 509192 432960
rect 509226 432926 509292 432960
rect 509326 432926 509392 432960
rect 509426 432926 510180 432960
rect 510214 432926 510280 432960
rect 510314 432926 510380 432960
rect 510414 432926 510480 432960
rect 510514 432926 510580 432960
rect 510614 432926 510680 432960
rect 510714 432926 511468 432960
rect 511502 432926 511568 432960
rect 511602 432926 511668 432960
rect 511702 432926 511768 432960
rect 511802 432926 511868 432960
rect 511902 432926 511968 432960
rect 512002 432926 512756 432960
rect 512790 432926 512856 432960
rect 512890 432926 512956 432960
rect 512990 432926 513056 432960
rect 513090 432926 513156 432960
rect 513190 432926 513256 432960
rect 513290 432926 513335 432960
rect 503709 432860 513335 432926
rect 503709 432826 503740 432860
rect 503774 432826 503840 432860
rect 503874 432826 503940 432860
rect 503974 432826 504040 432860
rect 504074 432826 504140 432860
rect 504174 432826 504240 432860
rect 504274 432826 505028 432860
rect 505062 432826 505128 432860
rect 505162 432826 505228 432860
rect 505262 432826 505328 432860
rect 505362 432826 505428 432860
rect 505462 432826 505528 432860
rect 505562 432826 506316 432860
rect 506350 432826 506416 432860
rect 506450 432826 506516 432860
rect 506550 432826 506616 432860
rect 506650 432826 506716 432860
rect 506750 432826 506816 432860
rect 506850 432826 507604 432860
rect 507638 432826 507704 432860
rect 507738 432826 507804 432860
rect 507838 432826 507904 432860
rect 507938 432826 508004 432860
rect 508038 432826 508104 432860
rect 508138 432826 508892 432860
rect 508926 432826 508992 432860
rect 509026 432826 509092 432860
rect 509126 432826 509192 432860
rect 509226 432826 509292 432860
rect 509326 432826 509392 432860
rect 509426 432826 510180 432860
rect 510214 432826 510280 432860
rect 510314 432826 510380 432860
rect 510414 432826 510480 432860
rect 510514 432826 510580 432860
rect 510614 432826 510680 432860
rect 510714 432826 511468 432860
rect 511502 432826 511568 432860
rect 511602 432826 511668 432860
rect 511702 432826 511768 432860
rect 511802 432826 511868 432860
rect 511902 432826 511968 432860
rect 512002 432826 512756 432860
rect 512790 432826 512856 432860
rect 512890 432826 512956 432860
rect 512990 432826 513056 432860
rect 513090 432826 513156 432860
rect 513190 432826 513256 432860
rect 513290 432826 513335 432860
rect 503709 432760 513335 432826
rect 503709 432726 503740 432760
rect 503774 432726 503840 432760
rect 503874 432726 503940 432760
rect 503974 432726 504040 432760
rect 504074 432726 504140 432760
rect 504174 432726 504240 432760
rect 504274 432726 505028 432760
rect 505062 432726 505128 432760
rect 505162 432726 505228 432760
rect 505262 432726 505328 432760
rect 505362 432726 505428 432760
rect 505462 432726 505528 432760
rect 505562 432726 506316 432760
rect 506350 432726 506416 432760
rect 506450 432726 506516 432760
rect 506550 432726 506616 432760
rect 506650 432726 506716 432760
rect 506750 432726 506816 432760
rect 506850 432726 507604 432760
rect 507638 432726 507704 432760
rect 507738 432726 507804 432760
rect 507838 432726 507904 432760
rect 507938 432726 508004 432760
rect 508038 432726 508104 432760
rect 508138 432726 508892 432760
rect 508926 432726 508992 432760
rect 509026 432726 509092 432760
rect 509126 432726 509192 432760
rect 509226 432726 509292 432760
rect 509326 432726 509392 432760
rect 509426 432726 510180 432760
rect 510214 432726 510280 432760
rect 510314 432726 510380 432760
rect 510414 432726 510480 432760
rect 510514 432726 510580 432760
rect 510614 432726 510680 432760
rect 510714 432726 511468 432760
rect 511502 432726 511568 432760
rect 511602 432726 511668 432760
rect 511702 432726 511768 432760
rect 511802 432726 511868 432760
rect 511902 432726 511968 432760
rect 512002 432726 512756 432760
rect 512790 432726 512856 432760
rect 512890 432726 512956 432760
rect 512990 432726 513056 432760
rect 513090 432726 513156 432760
rect 513190 432726 513256 432760
rect 513290 432726 513335 432760
rect 503709 432660 513335 432726
rect 503709 432626 503740 432660
rect 503774 432626 503840 432660
rect 503874 432626 503940 432660
rect 503974 432626 504040 432660
rect 504074 432626 504140 432660
rect 504174 432626 504240 432660
rect 504274 432626 505028 432660
rect 505062 432626 505128 432660
rect 505162 432626 505228 432660
rect 505262 432626 505328 432660
rect 505362 432626 505428 432660
rect 505462 432626 505528 432660
rect 505562 432626 506316 432660
rect 506350 432626 506416 432660
rect 506450 432626 506516 432660
rect 506550 432626 506616 432660
rect 506650 432626 506716 432660
rect 506750 432626 506816 432660
rect 506850 432626 507604 432660
rect 507638 432626 507704 432660
rect 507738 432626 507804 432660
rect 507838 432626 507904 432660
rect 507938 432626 508004 432660
rect 508038 432626 508104 432660
rect 508138 432626 508892 432660
rect 508926 432626 508992 432660
rect 509026 432626 509092 432660
rect 509126 432626 509192 432660
rect 509226 432626 509292 432660
rect 509326 432626 509392 432660
rect 509426 432626 510180 432660
rect 510214 432626 510280 432660
rect 510314 432626 510380 432660
rect 510414 432626 510480 432660
rect 510514 432626 510580 432660
rect 510614 432626 510680 432660
rect 510714 432626 511468 432660
rect 511502 432626 511568 432660
rect 511602 432626 511668 432660
rect 511702 432626 511768 432660
rect 511802 432626 511868 432660
rect 511902 432626 511968 432660
rect 512002 432626 512756 432660
rect 512790 432626 512856 432660
rect 512890 432626 512956 432660
rect 512990 432626 513056 432660
rect 513090 432626 513156 432660
rect 513190 432626 513256 432660
rect 513290 432626 513335 432660
rect 503709 432560 513335 432626
rect 503709 432526 503740 432560
rect 503774 432526 503840 432560
rect 503874 432526 503940 432560
rect 503974 432526 504040 432560
rect 504074 432526 504140 432560
rect 504174 432526 504240 432560
rect 504274 432526 505028 432560
rect 505062 432526 505128 432560
rect 505162 432526 505228 432560
rect 505262 432526 505328 432560
rect 505362 432526 505428 432560
rect 505462 432526 505528 432560
rect 505562 432526 506316 432560
rect 506350 432526 506416 432560
rect 506450 432526 506516 432560
rect 506550 432526 506616 432560
rect 506650 432526 506716 432560
rect 506750 432526 506816 432560
rect 506850 432526 507604 432560
rect 507638 432526 507704 432560
rect 507738 432526 507804 432560
rect 507838 432526 507904 432560
rect 507938 432526 508004 432560
rect 508038 432526 508104 432560
rect 508138 432526 508892 432560
rect 508926 432526 508992 432560
rect 509026 432526 509092 432560
rect 509126 432526 509192 432560
rect 509226 432526 509292 432560
rect 509326 432526 509392 432560
rect 509426 432526 510180 432560
rect 510214 432526 510280 432560
rect 510314 432526 510380 432560
rect 510414 432526 510480 432560
rect 510514 432526 510580 432560
rect 510614 432526 510680 432560
rect 510714 432526 511468 432560
rect 511502 432526 511568 432560
rect 511602 432526 511668 432560
rect 511702 432526 511768 432560
rect 511802 432526 511868 432560
rect 511902 432526 511968 432560
rect 512002 432526 512756 432560
rect 512790 432526 512856 432560
rect 512890 432526 512956 432560
rect 512990 432526 513056 432560
rect 513090 432526 513156 432560
rect 513190 432526 513256 432560
rect 513290 432526 513335 432560
rect 503709 432460 513335 432526
rect 503709 432426 503740 432460
rect 503774 432426 503840 432460
rect 503874 432426 503940 432460
rect 503974 432426 504040 432460
rect 504074 432426 504140 432460
rect 504174 432426 504240 432460
rect 504274 432426 505028 432460
rect 505062 432426 505128 432460
rect 505162 432426 505228 432460
rect 505262 432426 505328 432460
rect 505362 432426 505428 432460
rect 505462 432426 505528 432460
rect 505562 432426 506316 432460
rect 506350 432426 506416 432460
rect 506450 432426 506516 432460
rect 506550 432426 506616 432460
rect 506650 432426 506716 432460
rect 506750 432426 506816 432460
rect 506850 432426 507604 432460
rect 507638 432426 507704 432460
rect 507738 432426 507804 432460
rect 507838 432426 507904 432460
rect 507938 432426 508004 432460
rect 508038 432426 508104 432460
rect 508138 432426 508892 432460
rect 508926 432426 508992 432460
rect 509026 432426 509092 432460
rect 509126 432426 509192 432460
rect 509226 432426 509292 432460
rect 509326 432426 509392 432460
rect 509426 432426 510180 432460
rect 510214 432426 510280 432460
rect 510314 432426 510380 432460
rect 510414 432426 510480 432460
rect 510514 432426 510580 432460
rect 510614 432426 510680 432460
rect 510714 432426 511468 432460
rect 511502 432426 511568 432460
rect 511602 432426 511668 432460
rect 511702 432426 511768 432460
rect 511802 432426 511868 432460
rect 511902 432426 511968 432460
rect 512002 432426 512756 432460
rect 512790 432426 512856 432460
rect 512890 432426 512956 432460
rect 512990 432426 513056 432460
rect 513090 432426 513156 432460
rect 513190 432426 513256 432460
rect 513290 432426 513335 432460
rect 503709 432381 513335 432426
rect 527604 437540 528664 437580
rect 527604 437440 527638 437540
rect 527738 437440 527862 437540
rect 527962 437440 528086 437540
rect 528186 437440 528310 437540
rect 528410 437440 528534 437540
rect 528634 437440 528664 437540
rect 527604 437316 528664 437440
rect 527604 437216 527638 437316
rect 527738 437216 527862 437316
rect 527962 437216 528086 437316
rect 528186 437216 528310 437316
rect 528410 437216 528534 437316
rect 528634 437216 528664 437316
rect 527604 437092 528664 437216
rect 527604 436992 527638 437092
rect 527738 436992 527862 437092
rect 527962 436992 528086 437092
rect 528186 436992 528310 437092
rect 528410 436992 528534 437092
rect 528634 436992 528664 437092
rect 527604 436868 528664 436992
rect 527604 436768 527638 436868
rect 527738 436768 527862 436868
rect 527962 436768 528086 436868
rect 528186 436768 528310 436868
rect 528410 436768 528534 436868
rect 528634 436768 528664 436868
rect 527604 436644 528664 436768
rect 527604 436544 527638 436644
rect 527738 436544 527862 436644
rect 527962 436544 528086 436644
rect 528186 436544 528310 436644
rect 528410 436544 528534 436644
rect 528634 436544 528664 436644
rect 527604 436420 528664 436544
rect 527604 436320 527638 436420
rect 527738 436320 527862 436420
rect 527962 436320 528086 436420
rect 528186 436320 528310 436420
rect 528410 436320 528534 436420
rect 528634 436320 528664 436420
rect 527604 436196 528664 436320
rect 527604 436096 527638 436196
rect 527738 436096 527862 436196
rect 527962 436096 528086 436196
rect 528186 436096 528310 436196
rect 528410 436096 528534 436196
rect 528634 436096 528664 436196
rect 527604 435972 528664 436096
rect 527604 435872 527638 435972
rect 527738 435872 527862 435972
rect 527962 435872 528086 435972
rect 528186 435872 528310 435972
rect 528410 435872 528534 435972
rect 528634 435872 528664 435972
rect 527604 435748 528664 435872
rect 527604 435648 527638 435748
rect 527738 435648 527862 435748
rect 527962 435648 528086 435748
rect 528186 435648 528310 435748
rect 528410 435648 528534 435748
rect 528634 435648 528664 435748
rect 527604 435524 528664 435648
rect 527604 435424 527638 435524
rect 527738 435424 527862 435524
rect 527962 435424 528086 435524
rect 528186 435424 528310 435524
rect 528410 435424 528534 435524
rect 528634 435424 528664 435524
rect 527604 435300 528664 435424
rect 527604 435200 527638 435300
rect 527738 435200 527862 435300
rect 527962 435200 528086 435300
rect 528186 435200 528310 435300
rect 528410 435200 528534 435300
rect 528634 435200 528664 435300
rect 527604 435076 528664 435200
rect 527604 434976 527638 435076
rect 527738 434976 527862 435076
rect 527962 434976 528086 435076
rect 528186 434976 528310 435076
rect 528410 434976 528534 435076
rect 528634 434976 528664 435076
rect 527604 434852 528664 434976
rect 527604 434752 527638 434852
rect 527738 434752 527862 434852
rect 527962 434752 528086 434852
rect 528186 434752 528310 434852
rect 528410 434752 528534 434852
rect 528634 434752 528664 434852
rect 527604 434628 528664 434752
rect 527604 434528 527638 434628
rect 527738 434528 527862 434628
rect 527962 434528 528086 434628
rect 528186 434528 528310 434628
rect 528410 434528 528534 434628
rect 528634 434528 528664 434628
rect 527604 434404 528664 434528
rect 527604 434304 527638 434404
rect 527738 434304 527862 434404
rect 527962 434304 528086 434404
rect 528186 434304 528310 434404
rect 528410 434304 528534 434404
rect 528634 434304 528664 434404
rect 527604 434180 528664 434304
rect 527604 434080 527638 434180
rect 527738 434080 527862 434180
rect 527962 434080 528086 434180
rect 528186 434080 528310 434180
rect 528410 434080 528534 434180
rect 528634 434080 528664 434180
rect 527604 433956 528664 434080
rect 527604 433856 527638 433956
rect 527738 433856 527862 433956
rect 527962 433856 528086 433956
rect 528186 433856 528310 433956
rect 528410 433856 528534 433956
rect 528634 433856 528664 433956
rect 527604 433732 528664 433856
rect 527604 433632 527638 433732
rect 527738 433632 527862 433732
rect 527962 433632 528086 433732
rect 528186 433632 528310 433732
rect 528410 433632 528534 433732
rect 528634 433632 528664 433732
rect 527604 433508 528664 433632
rect 527604 433408 527638 433508
rect 527738 433408 527862 433508
rect 527962 433408 528086 433508
rect 528186 433408 528310 433508
rect 528410 433408 528534 433508
rect 528634 433408 528664 433508
rect 527604 433284 528664 433408
rect 527604 433184 527638 433284
rect 527738 433184 527862 433284
rect 527962 433184 528086 433284
rect 528186 433184 528310 433284
rect 528410 433184 528534 433284
rect 528634 433184 528664 433284
rect 527604 433060 528664 433184
rect 527604 432960 527638 433060
rect 527738 432960 527862 433060
rect 527962 432960 528086 433060
rect 528186 432960 528310 433060
rect 528410 432960 528534 433060
rect 528634 432960 528664 433060
rect 527604 432836 528664 432960
rect 527604 432736 527638 432836
rect 527738 432736 527862 432836
rect 527962 432736 528086 432836
rect 528186 432736 528310 432836
rect 528410 432736 528534 432836
rect 528634 432736 528664 432836
rect 527604 432612 528664 432736
rect 527604 432512 527638 432612
rect 527738 432512 527862 432612
rect 527962 432512 528086 432612
rect 528186 432512 528310 432612
rect 528410 432512 528534 432612
rect 528634 432512 528664 432612
rect 527604 432388 528664 432512
rect 500384 432164 501444 432288
rect 500384 432064 500418 432164
rect 500518 432064 500642 432164
rect 500742 432064 500866 432164
rect 500966 432064 501090 432164
rect 501190 432064 501314 432164
rect 501414 432064 501444 432164
rect 500384 431940 501444 432064
rect 500384 431840 500418 431940
rect 500518 431840 500642 431940
rect 500742 431840 500866 431940
rect 500966 431840 501090 431940
rect 501190 431840 501314 431940
rect 501414 431840 501444 431940
rect 500384 431716 501444 431840
rect 500384 431616 500418 431716
rect 500518 431616 500642 431716
rect 500742 431616 500866 431716
rect 500966 431616 501090 431716
rect 501190 431616 501314 431716
rect 501414 431616 501444 431716
rect 500384 431492 501444 431616
rect 500384 431392 500418 431492
rect 500518 431392 500642 431492
rect 500742 431392 500866 431492
rect 500966 431392 501090 431492
rect 501190 431392 501314 431492
rect 501414 431392 501444 431492
rect 500384 431268 501444 431392
rect 500384 431168 500418 431268
rect 500518 431168 500642 431268
rect 500742 431168 500866 431268
rect 500966 431168 501090 431268
rect 501190 431168 501314 431268
rect 501414 431168 501444 431268
rect 500384 431044 501444 431168
rect 527604 432288 527638 432388
rect 527738 432288 527862 432388
rect 527962 432288 528086 432388
rect 528186 432288 528310 432388
rect 528410 432288 528534 432388
rect 528634 432288 528664 432388
rect 527604 432164 528664 432288
rect 527604 432064 527638 432164
rect 527738 432064 527862 432164
rect 527962 432064 528086 432164
rect 528186 432064 528310 432164
rect 528410 432064 528534 432164
rect 528634 432064 528664 432164
rect 527604 431940 528664 432064
rect 527604 431840 527638 431940
rect 527738 431840 527862 431940
rect 527962 431840 528086 431940
rect 528186 431840 528310 431940
rect 528410 431840 528534 431940
rect 528634 431840 528664 431940
rect 527604 431716 528664 431840
rect 527604 431616 527638 431716
rect 527738 431616 527862 431716
rect 527962 431616 528086 431716
rect 528186 431616 528310 431716
rect 528410 431616 528534 431716
rect 528634 431616 528664 431716
rect 527604 431492 528664 431616
rect 527604 431392 527638 431492
rect 527738 431392 527862 431492
rect 527962 431392 528086 431492
rect 528186 431392 528310 431492
rect 528410 431392 528534 431492
rect 528634 431392 528664 431492
rect 527604 431268 528664 431392
rect 527604 431168 527638 431268
rect 527738 431168 527862 431268
rect 527962 431168 528086 431268
rect 528186 431168 528310 431268
rect 528410 431168 528534 431268
rect 528634 431168 528664 431268
rect 500384 430944 500418 431044
rect 500518 430944 500642 431044
rect 500742 430944 500866 431044
rect 500966 430944 501090 431044
rect 501190 430944 501314 431044
rect 501414 430944 501444 431044
rect 500384 430920 501444 430944
rect 503900 431026 510526 431056
rect 503900 430926 503920 431026
rect 504020 430926 504144 431026
rect 504244 430926 504368 431026
rect 504468 430926 504592 431026
rect 504692 430926 504816 431026
rect 504916 430926 505040 431026
rect 505140 430926 505264 431026
rect 505364 430926 505488 431026
rect 505588 430926 505712 431026
rect 505812 430926 505936 431026
rect 506036 430926 506160 431026
rect 506260 430926 506384 431026
rect 506484 430926 506608 431026
rect 506708 430926 506832 431026
rect 506932 430926 507056 431026
rect 507156 430926 507280 431026
rect 507380 430926 507504 431026
rect 507604 430926 507728 431026
rect 507828 430926 507952 431026
rect 508052 430926 508176 431026
rect 508276 430926 508400 431026
rect 508500 430926 508624 431026
rect 508724 430926 508848 431026
rect 508948 430926 509072 431026
rect 509172 430926 509296 431026
rect 509396 430926 509520 431026
rect 509620 430926 509744 431026
rect 509844 430926 509968 431026
rect 510068 430926 510192 431026
rect 510292 430926 510416 431026
rect 510516 430926 510526 431026
rect 503900 430802 510526 430926
rect 503900 430702 503920 430802
rect 504020 430702 504144 430802
rect 504244 430702 504368 430802
rect 504468 430702 504592 430802
rect 504692 430702 504816 430802
rect 504916 430702 505040 430802
rect 505140 430702 505264 430802
rect 505364 430702 505488 430802
rect 505588 430702 505712 430802
rect 505812 430702 505936 430802
rect 506036 430702 506160 430802
rect 506260 430702 506384 430802
rect 506484 430702 506608 430802
rect 506708 430702 506832 430802
rect 506932 430702 507056 430802
rect 507156 430702 507280 430802
rect 507380 430702 507504 430802
rect 507604 430702 507728 430802
rect 507828 430702 507952 430802
rect 508052 430702 508176 430802
rect 508276 430702 508400 430802
rect 508500 430702 508624 430802
rect 508724 430702 508848 430802
rect 508948 430702 509072 430802
rect 509172 430702 509296 430802
rect 509396 430702 509520 430802
rect 509620 430702 509744 430802
rect 509844 430702 509968 430802
rect 510068 430702 510192 430802
rect 510292 430702 510416 430802
rect 510516 430702 510526 430802
rect 503900 430578 510526 430702
rect 503900 430478 503920 430578
rect 504020 430478 504144 430578
rect 504244 430478 504368 430578
rect 504468 430478 504592 430578
rect 504692 430478 504816 430578
rect 504916 430478 505040 430578
rect 505140 430478 505264 430578
rect 505364 430478 505488 430578
rect 505588 430478 505712 430578
rect 505812 430478 505936 430578
rect 506036 430478 506160 430578
rect 506260 430478 506384 430578
rect 506484 430478 506608 430578
rect 506708 430478 506832 430578
rect 506932 430478 507056 430578
rect 507156 430478 507280 430578
rect 507380 430478 507504 430578
rect 507604 430478 507728 430578
rect 507828 430478 507952 430578
rect 508052 430478 508176 430578
rect 508276 430478 508400 430578
rect 508500 430478 508624 430578
rect 508724 430478 508848 430578
rect 508948 430478 509072 430578
rect 509172 430478 509296 430578
rect 509396 430478 509520 430578
rect 509620 430478 509744 430578
rect 509844 430478 509968 430578
rect 510068 430478 510192 430578
rect 510292 430478 510416 430578
rect 510516 430478 510526 430578
rect 503900 430354 510526 430478
rect 503900 430254 503920 430354
rect 504020 430254 504144 430354
rect 504244 430254 504368 430354
rect 504468 430254 504592 430354
rect 504692 430254 504816 430354
rect 504916 430254 505040 430354
rect 505140 430254 505264 430354
rect 505364 430254 505488 430354
rect 505588 430254 505712 430354
rect 505812 430254 505936 430354
rect 506036 430254 506160 430354
rect 506260 430254 506384 430354
rect 506484 430254 506608 430354
rect 506708 430254 506832 430354
rect 506932 430254 507056 430354
rect 507156 430254 507280 430354
rect 507380 430254 507504 430354
rect 507604 430254 507728 430354
rect 507828 430254 507952 430354
rect 508052 430254 508176 430354
rect 508276 430254 508400 430354
rect 508500 430254 508624 430354
rect 508724 430254 508848 430354
rect 508948 430254 509072 430354
rect 509172 430254 509296 430354
rect 509396 430254 509520 430354
rect 509620 430254 509744 430354
rect 509844 430254 509968 430354
rect 510068 430254 510192 430354
rect 510292 430254 510416 430354
rect 510516 430254 510526 430354
rect 503900 430130 510526 430254
rect 503900 430030 503920 430130
rect 504020 430030 504144 430130
rect 504244 430030 504368 430130
rect 504468 430030 504592 430130
rect 504692 430030 504816 430130
rect 504916 430030 505040 430130
rect 505140 430030 505264 430130
rect 505364 430030 505488 430130
rect 505588 430030 505712 430130
rect 505812 430030 505936 430130
rect 506036 430030 506160 430130
rect 506260 430030 506384 430130
rect 506484 430030 506608 430130
rect 506708 430030 506832 430130
rect 506932 430030 507056 430130
rect 507156 430030 507280 430130
rect 507380 430030 507504 430130
rect 507604 430030 507728 430130
rect 507828 430030 507952 430130
rect 508052 430030 508176 430130
rect 508276 430030 508400 430130
rect 508500 430030 508624 430130
rect 508724 430030 508848 430130
rect 508948 430030 509072 430130
rect 509172 430030 509296 430130
rect 509396 430030 509520 430130
rect 509620 430030 509744 430130
rect 509844 430030 509968 430130
rect 510068 430030 510192 430130
rect 510292 430030 510416 430130
rect 510516 430030 510526 430130
rect 503900 429998 510526 430030
rect 517280 431026 523940 431056
rect 517280 430926 517320 431026
rect 517420 430926 517544 431026
rect 517644 430926 517768 431026
rect 517868 430926 517992 431026
rect 518092 430926 518216 431026
rect 518316 430926 518440 431026
rect 518540 430926 518664 431026
rect 518764 430926 518888 431026
rect 518988 430926 519112 431026
rect 519212 430926 519336 431026
rect 519436 430926 519560 431026
rect 519660 430926 519784 431026
rect 519884 430926 520008 431026
rect 520108 430926 520232 431026
rect 520332 430926 520456 431026
rect 520556 430926 520680 431026
rect 520780 430926 520904 431026
rect 521004 430926 521128 431026
rect 521228 430926 521352 431026
rect 521452 430926 521576 431026
rect 521676 430926 521800 431026
rect 521900 430926 522024 431026
rect 522124 430926 522248 431026
rect 522348 430926 522472 431026
rect 522572 430926 522696 431026
rect 522796 430926 522920 431026
rect 523020 430926 523144 431026
rect 523244 430926 523368 431026
rect 523468 430926 523592 431026
rect 523692 430926 523816 431026
rect 523916 430926 523940 431026
rect 517280 430802 523940 430926
rect 527604 431044 528664 431168
rect 527604 430944 527638 431044
rect 527738 430944 527862 431044
rect 527962 430944 528086 431044
rect 528186 430944 528310 431044
rect 528410 430944 528534 431044
rect 528634 430944 528664 431044
rect 527604 430920 528664 430944
rect 517280 430702 517320 430802
rect 517420 430702 517544 430802
rect 517644 430702 517768 430802
rect 517868 430702 517992 430802
rect 518092 430702 518216 430802
rect 518316 430702 518440 430802
rect 518540 430702 518664 430802
rect 518764 430702 518888 430802
rect 518988 430702 519112 430802
rect 519212 430702 519336 430802
rect 519436 430702 519560 430802
rect 519660 430702 519784 430802
rect 519884 430702 520008 430802
rect 520108 430702 520232 430802
rect 520332 430702 520456 430802
rect 520556 430702 520680 430802
rect 520780 430702 520904 430802
rect 521004 430702 521128 430802
rect 521228 430702 521352 430802
rect 521452 430702 521576 430802
rect 521676 430702 521800 430802
rect 521900 430702 522024 430802
rect 522124 430702 522248 430802
rect 522348 430702 522472 430802
rect 522572 430702 522696 430802
rect 522796 430702 522920 430802
rect 523020 430702 523144 430802
rect 523244 430702 523368 430802
rect 523468 430702 523592 430802
rect 523692 430702 523816 430802
rect 523916 430702 523940 430802
rect 517280 430578 523940 430702
rect 517280 430478 517320 430578
rect 517420 430478 517544 430578
rect 517644 430478 517768 430578
rect 517868 430478 517992 430578
rect 518092 430478 518216 430578
rect 518316 430478 518440 430578
rect 518540 430478 518664 430578
rect 518764 430478 518888 430578
rect 518988 430478 519112 430578
rect 519212 430478 519336 430578
rect 519436 430478 519560 430578
rect 519660 430478 519784 430578
rect 519884 430478 520008 430578
rect 520108 430478 520232 430578
rect 520332 430478 520456 430578
rect 520556 430478 520680 430578
rect 520780 430478 520904 430578
rect 521004 430478 521128 430578
rect 521228 430478 521352 430578
rect 521452 430478 521576 430578
rect 521676 430478 521800 430578
rect 521900 430478 522024 430578
rect 522124 430478 522248 430578
rect 522348 430478 522472 430578
rect 522572 430478 522696 430578
rect 522796 430478 522920 430578
rect 523020 430478 523144 430578
rect 523244 430478 523368 430578
rect 523468 430478 523592 430578
rect 523692 430478 523816 430578
rect 523916 430478 523940 430578
rect 517280 430354 523940 430478
rect 517280 430254 517320 430354
rect 517420 430254 517544 430354
rect 517644 430254 517768 430354
rect 517868 430254 517992 430354
rect 518092 430254 518216 430354
rect 518316 430254 518440 430354
rect 518540 430254 518664 430354
rect 518764 430254 518888 430354
rect 518988 430254 519112 430354
rect 519212 430254 519336 430354
rect 519436 430254 519560 430354
rect 519660 430254 519784 430354
rect 519884 430254 520008 430354
rect 520108 430254 520232 430354
rect 520332 430254 520456 430354
rect 520556 430254 520680 430354
rect 520780 430254 520904 430354
rect 521004 430254 521128 430354
rect 521228 430254 521352 430354
rect 521452 430254 521576 430354
rect 521676 430254 521800 430354
rect 521900 430254 522024 430354
rect 522124 430254 522248 430354
rect 522348 430254 522472 430354
rect 522572 430254 522696 430354
rect 522796 430254 522920 430354
rect 523020 430254 523144 430354
rect 523244 430254 523368 430354
rect 523468 430254 523592 430354
rect 523692 430254 523816 430354
rect 523916 430254 523940 430354
rect 517280 430130 523940 430254
rect 517280 430030 517320 430130
rect 517420 430030 517544 430130
rect 517644 430030 517768 430130
rect 517868 430030 517992 430130
rect 518092 430030 518216 430130
rect 518316 430030 518440 430130
rect 518540 430030 518664 430130
rect 518764 430030 518888 430130
rect 518988 430030 519112 430130
rect 519212 430030 519336 430130
rect 519436 430030 519560 430130
rect 519660 430030 519784 430130
rect 519884 430030 520008 430130
rect 520108 430030 520232 430130
rect 520332 430030 520456 430130
rect 520556 430030 520680 430130
rect 520780 430030 520904 430130
rect 521004 430030 521128 430130
rect 521228 430030 521352 430130
rect 521452 430030 521576 430130
rect 521676 430030 521800 430130
rect 521900 430030 522024 430130
rect 522124 430030 522248 430130
rect 522348 430030 522472 430130
rect 522572 430030 522696 430130
rect 522796 430030 522920 430130
rect 523020 430030 523144 430130
rect 523244 430030 523368 430130
rect 523468 430030 523592 430130
rect 523692 430030 523816 430130
rect 523916 430030 523940 430130
rect 517280 429996 523940 430030
<< via1 >>
rect 562480 495662 562560 495742
rect 562640 495662 562720 495742
rect 562800 495662 562880 495742
rect 562960 495662 563040 495742
rect 563120 495662 563200 495742
rect 563280 495662 563360 495742
rect 563440 495662 563520 495742
rect 563600 495662 563680 495742
rect 563760 495662 563840 495742
rect 563920 495662 564000 495742
rect 564080 495662 564160 495742
rect 564240 495662 564320 495742
rect 564400 495662 564480 495742
rect 564560 495662 564640 495742
rect 564720 495662 564800 495742
rect 564880 495662 564960 495742
rect 565040 495662 565120 495742
rect 565200 495662 565280 495742
rect 565360 495662 565440 495742
rect 565520 495662 565600 495742
rect 565680 495662 565760 495742
rect 565840 495662 565920 495742
rect 566000 495662 566080 495742
rect 566160 495662 566240 495742
rect 566320 495662 566400 495742
rect 566480 495662 566560 495742
rect 566640 495662 566720 495742
rect 566800 495662 566880 495742
rect 566960 495662 567040 495742
rect 567120 495662 567200 495742
rect 567280 495662 567360 495742
rect 562480 495514 562560 495582
rect 562640 495514 562720 495582
rect 562800 495514 562880 495582
rect 562960 495514 563040 495582
rect 563120 495514 563200 495582
rect 563280 495514 563360 495582
rect 563440 495514 563520 495582
rect 563600 495514 563680 495582
rect 563760 495514 563840 495582
rect 563920 495514 564000 495582
rect 564080 495514 564160 495582
rect 564240 495514 564320 495582
rect 564400 495514 564480 495582
rect 564560 495514 564640 495582
rect 564720 495514 564800 495582
rect 564880 495514 564960 495582
rect 565040 495514 565120 495582
rect 565200 495514 565280 495582
rect 565360 495514 565440 495582
rect 565520 495514 565600 495582
rect 565680 495514 565760 495582
rect 565840 495514 565920 495582
rect 566000 495514 566080 495582
rect 566160 495514 566240 495582
rect 566320 495514 566400 495582
rect 566480 495514 566560 495582
rect 566640 495514 566720 495582
rect 566800 495514 566880 495582
rect 566960 495514 567040 495582
rect 567120 495514 567200 495582
rect 567280 495514 567360 495582
rect 562480 495502 562560 495514
rect 562640 495502 562720 495514
rect 562800 495502 562880 495514
rect 562960 495502 563040 495514
rect 563120 495502 563200 495514
rect 563280 495502 563360 495514
rect 563440 495502 563520 495514
rect 563600 495502 563680 495514
rect 563760 495502 563840 495514
rect 563920 495502 564000 495514
rect 564080 495502 564160 495514
rect 564240 495502 564320 495514
rect 564400 495502 564480 495514
rect 564560 495502 564640 495514
rect 564720 495502 564800 495514
rect 564880 495502 564960 495514
rect 565040 495502 565120 495514
rect 565200 495502 565280 495514
rect 565360 495502 565440 495514
rect 565520 495502 565600 495514
rect 565680 495502 565760 495514
rect 565840 495502 565920 495514
rect 566000 495502 566080 495514
rect 566160 495502 566240 495514
rect 566320 495502 566400 495514
rect 566480 495502 566560 495514
rect 566640 495502 566720 495514
rect 566800 495502 566880 495514
rect 566960 495502 567040 495514
rect 567120 495502 567200 495514
rect 567280 495502 567360 495514
rect 572640 495662 572720 495742
rect 572800 495662 572880 495742
rect 572960 495662 573040 495742
rect 573120 495662 573200 495742
rect 573280 495662 573360 495742
rect 573440 495662 573520 495742
rect 573600 495662 573680 495742
rect 573760 495662 573840 495742
rect 573920 495662 574000 495742
rect 574080 495662 574160 495742
rect 574240 495662 574320 495742
rect 574400 495662 574480 495742
rect 574560 495662 574640 495742
rect 574720 495662 574800 495742
rect 574880 495662 574960 495742
rect 575040 495662 575120 495742
rect 575200 495662 575280 495742
rect 575360 495662 575440 495742
rect 575520 495662 575600 495742
rect 575680 495662 575760 495742
rect 575840 495662 575920 495742
rect 576000 495662 576080 495742
rect 576160 495662 576240 495742
rect 576320 495662 576400 495742
rect 576480 495662 576560 495742
rect 576640 495662 576720 495742
rect 576800 495662 576880 495742
rect 576960 495662 577040 495742
rect 577120 495662 577200 495742
rect 577280 495662 577360 495742
rect 577440 495662 577520 495742
rect 572640 495548 572720 495582
rect 572800 495548 572880 495582
rect 572960 495548 573040 495582
rect 573120 495548 573200 495582
rect 573280 495548 573360 495582
rect 573440 495548 573520 495582
rect 573600 495548 573680 495582
rect 573760 495548 573840 495582
rect 573920 495548 574000 495582
rect 574080 495548 574160 495582
rect 574240 495548 574320 495582
rect 574400 495548 574480 495582
rect 574560 495548 574640 495582
rect 574720 495548 574800 495582
rect 574880 495548 574960 495582
rect 575040 495548 575120 495582
rect 575200 495548 575280 495582
rect 575360 495548 575440 495582
rect 575520 495548 575600 495582
rect 575680 495548 575760 495582
rect 575840 495548 575920 495582
rect 576000 495548 576080 495582
rect 576160 495548 576240 495582
rect 576320 495548 576400 495582
rect 576480 495548 576560 495582
rect 576640 495548 576720 495582
rect 576800 495548 576880 495582
rect 576960 495548 577040 495582
rect 577120 495548 577200 495582
rect 577280 495548 577360 495582
rect 577440 495548 577520 495582
rect 572640 495514 572720 495548
rect 572800 495514 572880 495548
rect 572960 495514 573040 495548
rect 573120 495514 573200 495548
rect 573280 495514 573360 495548
rect 573440 495514 573520 495548
rect 573600 495514 573680 495548
rect 573760 495514 573840 495548
rect 573920 495514 574000 495548
rect 574080 495514 574160 495548
rect 574240 495514 574320 495548
rect 574400 495514 574480 495548
rect 574560 495514 574640 495548
rect 574720 495514 574800 495548
rect 574880 495514 574960 495548
rect 575040 495514 575120 495548
rect 575200 495514 575280 495548
rect 575360 495514 575440 495548
rect 575520 495514 575600 495548
rect 575680 495514 575760 495548
rect 575840 495514 575920 495548
rect 576000 495514 576080 495548
rect 576160 495514 576240 495548
rect 576320 495514 576400 495548
rect 576480 495514 576560 495548
rect 576640 495514 576720 495548
rect 576800 495514 576880 495548
rect 576960 495514 577040 495548
rect 577120 495514 577200 495548
rect 577280 495514 577360 495548
rect 577440 495514 577520 495548
rect 572640 495502 572720 495514
rect 572800 495502 572880 495514
rect 572960 495502 573040 495514
rect 573120 495502 573200 495514
rect 573280 495502 573360 495514
rect 573440 495502 573520 495514
rect 573600 495502 573680 495514
rect 573760 495502 573840 495514
rect 573920 495502 574000 495514
rect 574080 495502 574160 495514
rect 574240 495502 574320 495514
rect 574400 495502 574480 495514
rect 574560 495502 574640 495514
rect 574720 495502 574800 495514
rect 574880 495502 574960 495514
rect 575040 495502 575120 495514
rect 575200 495502 575280 495514
rect 575360 495502 575440 495514
rect 575520 495502 575600 495514
rect 575680 495502 575760 495514
rect 575840 495502 575920 495514
rect 576000 495502 576080 495514
rect 576160 495502 576240 495514
rect 576320 495502 576400 495514
rect 576480 495502 576560 495514
rect 576640 495502 576720 495514
rect 576800 495502 576880 495514
rect 576960 495502 577040 495514
rect 577120 495502 577200 495514
rect 577280 495502 577360 495514
rect 577440 495502 577520 495514
rect 562222 494161 562282 494221
rect 562342 494161 562402 494221
rect 562462 494161 562522 494221
rect 562582 494161 562642 494221
rect 562702 494161 562762 494221
rect 562822 494161 562882 494221
rect 562942 494161 563002 494221
rect 563062 494161 563122 494221
rect 563182 494161 563242 494221
rect 563302 494161 563362 494221
rect 563422 494161 563482 494221
rect 563542 494161 563602 494221
rect 563662 494161 563722 494221
rect 563782 494161 563842 494221
rect 563902 494161 563962 494221
rect 564022 494161 564082 494221
rect 564142 494161 564202 494221
rect 564262 494161 564322 494221
rect 564382 494161 564442 494221
rect 564502 494161 564562 494221
rect 564622 494161 564682 494221
rect 564742 494161 564802 494221
rect 564862 494161 564922 494221
rect 564982 494161 565042 494221
rect 565102 494161 565162 494221
rect 565222 494161 565282 494221
rect 565342 494161 565402 494221
rect 565462 494161 565522 494221
rect 565582 494161 565642 494221
rect 565702 494161 565762 494221
rect 565822 494161 565882 494221
rect 565942 494161 566002 494221
rect 566062 494161 566122 494221
rect 566182 494161 566242 494221
rect 566302 494161 566362 494221
rect 566422 494161 566482 494221
rect 566542 494161 566602 494221
rect 566662 494161 566722 494221
rect 566782 494161 566842 494221
rect 566902 494161 566962 494221
rect 567022 494161 567082 494221
rect 567142 494161 567202 494221
rect 567262 494161 567322 494221
rect 567382 494161 567442 494221
rect 567502 494161 567562 494221
rect 562222 494041 562282 494101
rect 562342 494041 562402 494101
rect 562462 494041 562522 494101
rect 562582 494041 562642 494101
rect 562702 494041 562762 494101
rect 562822 494041 562882 494101
rect 562942 494041 563002 494101
rect 563062 494041 563122 494101
rect 563182 494041 563242 494101
rect 563302 494041 563362 494101
rect 563422 494041 563482 494101
rect 563542 494041 563602 494101
rect 563662 494041 563722 494101
rect 563782 494041 563842 494101
rect 563902 494041 563962 494101
rect 564022 494041 564082 494101
rect 564142 494041 564202 494101
rect 564262 494041 564322 494101
rect 564382 494041 564442 494101
rect 564502 494041 564562 494101
rect 564622 494041 564682 494101
rect 564742 494041 564802 494101
rect 564862 494041 564922 494101
rect 564982 494041 565042 494101
rect 565102 494041 565162 494101
rect 565222 494041 565282 494101
rect 565342 494041 565402 494101
rect 565462 494041 565522 494101
rect 565582 494041 565642 494101
rect 565702 494041 565762 494101
rect 565822 494041 565882 494101
rect 565942 494041 566002 494101
rect 566062 494041 566122 494101
rect 566182 494041 566242 494101
rect 566302 494041 566362 494101
rect 566422 494041 566482 494101
rect 566542 494041 566602 494101
rect 566662 494041 566722 494101
rect 566782 494041 566842 494101
rect 566902 494041 566962 494101
rect 567022 494041 567082 494101
rect 567142 494041 567202 494101
rect 567262 494041 567322 494101
rect 567382 494041 567442 494101
rect 567502 494041 567562 494101
rect 572332 494176 572392 494236
rect 572452 494176 572512 494236
rect 572572 494176 572632 494236
rect 572692 494176 572752 494236
rect 572812 494176 572872 494236
rect 572932 494176 572992 494236
rect 573052 494176 573112 494236
rect 573172 494176 573232 494236
rect 573292 494176 573352 494236
rect 573412 494176 573472 494236
rect 573532 494176 573592 494236
rect 573652 494176 573712 494236
rect 573772 494176 573832 494236
rect 573892 494176 573952 494236
rect 574012 494176 574072 494236
rect 574132 494176 574192 494236
rect 574252 494176 574312 494236
rect 574372 494176 574432 494236
rect 574492 494176 574552 494236
rect 574612 494176 574672 494236
rect 574732 494176 574792 494236
rect 574852 494176 574912 494236
rect 574972 494176 575032 494236
rect 575092 494176 575152 494236
rect 575212 494176 575272 494236
rect 575332 494176 575392 494236
rect 575452 494176 575512 494236
rect 575572 494176 575632 494236
rect 575692 494176 575752 494236
rect 575812 494176 575872 494236
rect 575932 494176 575992 494236
rect 576052 494176 576112 494236
rect 576172 494176 576232 494236
rect 576292 494176 576352 494236
rect 576412 494176 576472 494236
rect 576532 494176 576592 494236
rect 576652 494176 576712 494236
rect 576772 494176 576832 494236
rect 576892 494176 576952 494236
rect 577012 494176 577072 494236
rect 577132 494176 577192 494236
rect 577252 494176 577312 494236
rect 577372 494176 577432 494236
rect 577492 494176 577552 494236
rect 577612 494176 577672 494236
rect 572332 494056 572392 494116
rect 572452 494056 572512 494116
rect 572572 494056 572632 494116
rect 572692 494056 572752 494116
rect 572812 494056 572872 494116
rect 572932 494056 572992 494116
rect 573052 494056 573112 494116
rect 573172 494056 573232 494116
rect 573292 494056 573352 494116
rect 573412 494056 573472 494116
rect 573532 494056 573592 494116
rect 573652 494056 573712 494116
rect 573772 494056 573832 494116
rect 573892 494056 573952 494116
rect 574012 494056 574072 494116
rect 574132 494056 574192 494116
rect 574252 494056 574312 494116
rect 574372 494056 574432 494116
rect 574492 494056 574552 494116
rect 574612 494056 574672 494116
rect 574732 494056 574792 494116
rect 574852 494056 574912 494116
rect 574972 494056 575032 494116
rect 575092 494056 575152 494116
rect 575212 494056 575272 494116
rect 575332 494056 575392 494116
rect 575452 494056 575512 494116
rect 575572 494056 575632 494116
rect 575692 494056 575752 494116
rect 575812 494056 575872 494116
rect 575932 494056 575992 494116
rect 576052 494056 576112 494116
rect 576172 494056 576232 494116
rect 576292 494056 576352 494116
rect 576412 494056 576472 494116
rect 576532 494056 576592 494116
rect 576652 494056 576712 494116
rect 576772 494056 576832 494116
rect 576892 494056 576952 494116
rect 577012 494056 577072 494116
rect 577132 494056 577192 494116
rect 577252 494056 577312 494116
rect 577372 494056 577432 494116
rect 577492 494056 577552 494116
rect 577612 494056 577672 494116
rect 503920 475206 504020 475306
rect 504144 475206 504244 475306
rect 504368 475206 504468 475306
rect 504592 475206 504692 475306
rect 504816 475206 504916 475306
rect 505040 475206 505140 475306
rect 505264 475206 505364 475306
rect 505488 475206 505588 475306
rect 505712 475206 505812 475306
rect 505936 475206 506036 475306
rect 506160 475206 506260 475306
rect 506384 475206 506484 475306
rect 506608 475206 506708 475306
rect 506832 475206 506932 475306
rect 507056 475206 507156 475306
rect 507280 475206 507380 475306
rect 507504 475206 507604 475306
rect 507728 475206 507828 475306
rect 507952 475206 508052 475306
rect 508176 475206 508276 475306
rect 508400 475206 508500 475306
rect 508624 475206 508724 475306
rect 508848 475206 508948 475306
rect 509072 475206 509172 475306
rect 509296 475206 509396 475306
rect 509520 475206 509620 475306
rect 509744 475206 509844 475306
rect 509968 475206 510068 475306
rect 510192 475206 510292 475306
rect 510416 475206 510516 475306
rect 503920 474982 504020 475082
rect 504144 474982 504244 475082
rect 504368 474982 504468 475082
rect 504592 474982 504692 475082
rect 504816 474982 504916 475082
rect 505040 474982 505140 475082
rect 505264 474982 505364 475082
rect 505488 474982 505588 475082
rect 505712 474982 505812 475082
rect 505936 474982 506036 475082
rect 506160 474982 506260 475082
rect 506384 474982 506484 475082
rect 506608 474982 506708 475082
rect 506832 474982 506932 475082
rect 507056 474982 507156 475082
rect 507280 474982 507380 475082
rect 507504 474982 507604 475082
rect 507728 474982 507828 475082
rect 507952 474982 508052 475082
rect 508176 474982 508276 475082
rect 508400 474982 508500 475082
rect 508624 474982 508724 475082
rect 508848 474982 508948 475082
rect 509072 474982 509172 475082
rect 509296 474982 509396 475082
rect 509520 474982 509620 475082
rect 509744 474982 509844 475082
rect 509968 474982 510068 475082
rect 510192 474982 510292 475082
rect 510416 474982 510516 475082
rect 503920 474758 504020 474858
rect 504144 474758 504244 474858
rect 504368 474758 504468 474858
rect 504592 474758 504692 474858
rect 504816 474758 504916 474858
rect 505040 474758 505140 474858
rect 505264 474758 505364 474858
rect 505488 474758 505588 474858
rect 505712 474758 505812 474858
rect 505936 474758 506036 474858
rect 506160 474758 506260 474858
rect 506384 474758 506484 474858
rect 506608 474758 506708 474858
rect 506832 474758 506932 474858
rect 507056 474758 507156 474858
rect 507280 474758 507380 474858
rect 507504 474758 507604 474858
rect 507728 474758 507828 474858
rect 507952 474758 508052 474858
rect 508176 474758 508276 474858
rect 508400 474758 508500 474858
rect 508624 474758 508724 474858
rect 508848 474758 508948 474858
rect 509072 474758 509172 474858
rect 509296 474758 509396 474858
rect 509520 474758 509620 474858
rect 509744 474758 509844 474858
rect 509968 474758 510068 474858
rect 510192 474758 510292 474858
rect 510416 474758 510516 474858
rect 503920 474534 504020 474634
rect 504144 474534 504244 474634
rect 504368 474534 504468 474634
rect 504592 474534 504692 474634
rect 504816 474534 504916 474634
rect 505040 474534 505140 474634
rect 505264 474534 505364 474634
rect 505488 474534 505588 474634
rect 505712 474534 505812 474634
rect 505936 474534 506036 474634
rect 506160 474534 506260 474634
rect 506384 474534 506484 474634
rect 506608 474534 506708 474634
rect 506832 474534 506932 474634
rect 507056 474534 507156 474634
rect 507280 474534 507380 474634
rect 507504 474534 507604 474634
rect 507728 474534 507828 474634
rect 507952 474534 508052 474634
rect 508176 474534 508276 474634
rect 508400 474534 508500 474634
rect 508624 474534 508724 474634
rect 508848 474534 508948 474634
rect 509072 474534 509172 474634
rect 509296 474534 509396 474634
rect 509520 474534 509620 474634
rect 509744 474534 509844 474634
rect 509968 474534 510068 474634
rect 510192 474534 510292 474634
rect 510416 474534 510516 474634
rect 500398 474180 500498 474280
rect 500622 474180 500722 474280
rect 500846 474180 500946 474280
rect 501070 474180 501170 474280
rect 501294 474180 501394 474280
rect 503920 474310 504020 474410
rect 504144 474310 504244 474410
rect 504368 474310 504468 474410
rect 504592 474310 504692 474410
rect 504816 474310 504916 474410
rect 505040 474310 505140 474410
rect 505264 474310 505364 474410
rect 505488 474310 505588 474410
rect 505712 474310 505812 474410
rect 505936 474310 506036 474410
rect 506160 474310 506260 474410
rect 506384 474310 506484 474410
rect 506608 474310 506708 474410
rect 506832 474310 506932 474410
rect 507056 474310 507156 474410
rect 507280 474310 507380 474410
rect 507504 474310 507604 474410
rect 507728 474310 507828 474410
rect 507952 474310 508052 474410
rect 508176 474310 508276 474410
rect 508400 474310 508500 474410
rect 508624 474310 508724 474410
rect 508848 474310 508948 474410
rect 509072 474310 509172 474410
rect 509296 474310 509396 474410
rect 509520 474310 509620 474410
rect 509744 474310 509844 474410
rect 509968 474310 510068 474410
rect 510192 474310 510292 474410
rect 510416 474310 510516 474410
rect 517320 475206 517420 475306
rect 517544 475206 517644 475306
rect 517768 475206 517868 475306
rect 517992 475206 518092 475306
rect 518216 475206 518316 475306
rect 518440 475206 518540 475306
rect 518664 475206 518764 475306
rect 518888 475206 518988 475306
rect 519112 475206 519212 475306
rect 519336 475206 519436 475306
rect 519560 475206 519660 475306
rect 519784 475206 519884 475306
rect 520008 475206 520108 475306
rect 520232 475206 520332 475306
rect 520456 475206 520556 475306
rect 520680 475206 520780 475306
rect 520904 475206 521004 475306
rect 521128 475206 521228 475306
rect 521352 475206 521452 475306
rect 521576 475206 521676 475306
rect 521800 475206 521900 475306
rect 522024 475206 522124 475306
rect 522248 475206 522348 475306
rect 522472 475206 522572 475306
rect 522696 475206 522796 475306
rect 522920 475206 523020 475306
rect 523144 475206 523244 475306
rect 523368 475206 523468 475306
rect 523592 475206 523692 475306
rect 523816 475206 523916 475306
rect 517320 474982 517420 475082
rect 517544 474982 517644 475082
rect 517768 474982 517868 475082
rect 517992 474982 518092 475082
rect 518216 474982 518316 475082
rect 518440 474982 518540 475082
rect 518664 474982 518764 475082
rect 518888 474982 518988 475082
rect 519112 474982 519212 475082
rect 519336 474982 519436 475082
rect 519560 474982 519660 475082
rect 519784 474982 519884 475082
rect 520008 474982 520108 475082
rect 520232 474982 520332 475082
rect 520456 474982 520556 475082
rect 520680 474982 520780 475082
rect 520904 474982 521004 475082
rect 521128 474982 521228 475082
rect 521352 474982 521452 475082
rect 521576 474982 521676 475082
rect 521800 474982 521900 475082
rect 522024 474982 522124 475082
rect 522248 474982 522348 475082
rect 522472 474982 522572 475082
rect 522696 474982 522796 475082
rect 522920 474982 523020 475082
rect 523144 474982 523244 475082
rect 523368 474982 523468 475082
rect 523592 474982 523692 475082
rect 523816 474982 523916 475082
rect 517320 474758 517420 474858
rect 517544 474758 517644 474858
rect 517768 474758 517868 474858
rect 517992 474758 518092 474858
rect 518216 474758 518316 474858
rect 518440 474758 518540 474858
rect 518664 474758 518764 474858
rect 518888 474758 518988 474858
rect 519112 474758 519212 474858
rect 519336 474758 519436 474858
rect 519560 474758 519660 474858
rect 519784 474758 519884 474858
rect 520008 474758 520108 474858
rect 520232 474758 520332 474858
rect 520456 474758 520556 474858
rect 520680 474758 520780 474858
rect 520904 474758 521004 474858
rect 521128 474758 521228 474858
rect 521352 474758 521452 474858
rect 521576 474758 521676 474858
rect 521800 474758 521900 474858
rect 522024 474758 522124 474858
rect 522248 474758 522348 474858
rect 522472 474758 522572 474858
rect 522696 474758 522796 474858
rect 522920 474758 523020 474858
rect 523144 474758 523244 474858
rect 523368 474758 523468 474858
rect 523592 474758 523692 474858
rect 523816 474758 523916 474858
rect 517320 474534 517420 474634
rect 517544 474534 517644 474634
rect 517768 474534 517868 474634
rect 517992 474534 518092 474634
rect 518216 474534 518316 474634
rect 518440 474534 518540 474634
rect 518664 474534 518764 474634
rect 518888 474534 518988 474634
rect 519112 474534 519212 474634
rect 519336 474534 519436 474634
rect 519560 474534 519660 474634
rect 519784 474534 519884 474634
rect 520008 474534 520108 474634
rect 520232 474534 520332 474634
rect 520456 474534 520556 474634
rect 520680 474534 520780 474634
rect 520904 474534 521004 474634
rect 521128 474534 521228 474634
rect 521352 474534 521452 474634
rect 521576 474534 521676 474634
rect 521800 474534 521900 474634
rect 522024 474534 522124 474634
rect 522248 474534 522348 474634
rect 522472 474534 522572 474634
rect 522696 474534 522796 474634
rect 522920 474534 523020 474634
rect 523144 474534 523244 474634
rect 523368 474534 523468 474634
rect 523592 474534 523692 474634
rect 523816 474534 523916 474634
rect 517320 474310 517420 474410
rect 517544 474310 517644 474410
rect 517768 474310 517868 474410
rect 517992 474310 518092 474410
rect 518216 474310 518316 474410
rect 518440 474310 518540 474410
rect 518664 474310 518764 474410
rect 518888 474310 518988 474410
rect 519112 474310 519212 474410
rect 519336 474310 519436 474410
rect 519560 474310 519660 474410
rect 519784 474310 519884 474410
rect 520008 474310 520108 474410
rect 520232 474310 520332 474410
rect 520456 474310 520556 474410
rect 520680 474310 520780 474410
rect 520904 474310 521004 474410
rect 521128 474310 521228 474410
rect 521352 474310 521452 474410
rect 521576 474310 521676 474410
rect 521800 474310 521900 474410
rect 522024 474310 522124 474410
rect 522248 474310 522348 474410
rect 522472 474310 522572 474410
rect 522696 474310 522796 474410
rect 522920 474310 523020 474410
rect 523144 474310 523244 474410
rect 523368 474310 523468 474410
rect 523592 474310 523692 474410
rect 523816 474310 523916 474410
rect 500398 473956 500498 474056
rect 500622 473956 500722 474056
rect 500846 473956 500946 474056
rect 501070 473956 501170 474056
rect 501294 473956 501394 474056
rect 500398 473732 500498 473832
rect 500622 473732 500722 473832
rect 500846 473732 500946 473832
rect 501070 473732 501170 473832
rect 501294 473732 501394 473832
rect 500398 473508 500498 473608
rect 500622 473508 500722 473608
rect 500846 473508 500946 473608
rect 501070 473508 501170 473608
rect 501294 473508 501394 473608
rect 500398 473284 500498 473384
rect 500622 473284 500722 473384
rect 500846 473284 500946 473384
rect 501070 473284 501170 473384
rect 501294 473284 501394 473384
rect 500398 473060 500498 473160
rect 500622 473060 500722 473160
rect 500846 473060 500946 473160
rect 501070 473060 501170 473160
rect 501294 473060 501394 473160
rect 500398 472836 500498 472936
rect 500622 472836 500722 472936
rect 500846 472836 500946 472936
rect 501070 472836 501170 472936
rect 501294 472836 501394 472936
rect 527618 474180 527718 474280
rect 527842 474180 527942 474280
rect 528066 474180 528166 474280
rect 528290 474180 528390 474280
rect 528514 474180 528614 474280
rect 527618 473956 527718 474056
rect 527842 473956 527942 474056
rect 528066 473956 528166 474056
rect 528290 473956 528390 474056
rect 528514 473956 528614 474056
rect 527618 473732 527718 473832
rect 527842 473732 527942 473832
rect 528066 473732 528166 473832
rect 528290 473732 528390 473832
rect 528514 473732 528614 473832
rect 527618 473508 527718 473608
rect 527842 473508 527942 473608
rect 528066 473508 528166 473608
rect 528290 473508 528390 473608
rect 528514 473508 528614 473608
rect 527618 473284 527718 473384
rect 527842 473284 527942 473384
rect 528066 473284 528166 473384
rect 528290 473284 528390 473384
rect 528514 473284 528614 473384
rect 527618 473060 527718 473160
rect 527842 473060 527942 473160
rect 528066 473060 528166 473160
rect 528290 473060 528390 473160
rect 528514 473060 528614 473160
rect 527618 472836 527718 472936
rect 527842 472836 527942 472936
rect 528066 472836 528166 472936
rect 528290 472836 528390 472936
rect 528514 472836 528614 472936
rect 500398 472612 500498 472712
rect 500622 472612 500722 472712
rect 500846 472612 500946 472712
rect 501070 472612 501170 472712
rect 501294 472612 501394 472712
rect 500398 472388 500498 472488
rect 500622 472388 500722 472488
rect 500846 472388 500946 472488
rect 501070 472388 501170 472488
rect 501294 472388 501394 472488
rect 527618 472612 527718 472712
rect 527842 472612 527942 472712
rect 528066 472612 528166 472712
rect 528290 472612 528390 472712
rect 528514 472612 528614 472712
rect 500398 472164 500498 472264
rect 500622 472164 500722 472264
rect 500846 472164 500946 472264
rect 501070 472164 501170 472264
rect 501294 472164 501394 472264
rect 506370 472264 506422 472316
rect 500398 471940 500498 472040
rect 500622 471940 500722 472040
rect 500846 471940 500946 472040
rect 501070 471940 501170 472040
rect 501294 471940 501394 472040
rect 500398 471716 500498 471816
rect 500622 471716 500722 471816
rect 500846 471716 500946 471816
rect 501070 471716 501170 471816
rect 501294 471716 501394 471816
rect 500398 471492 500498 471592
rect 500622 471492 500722 471592
rect 500846 471492 500946 471592
rect 501070 471492 501170 471592
rect 501294 471492 501394 471592
rect 500398 471268 500498 471368
rect 500622 471268 500722 471368
rect 500846 471268 500946 471368
rect 501070 471268 501170 471368
rect 501294 471268 501394 471368
rect 506164 471346 506216 471398
rect 500398 471044 500498 471144
rect 500622 471044 500722 471144
rect 500846 471044 500946 471144
rect 501070 471044 501170 471144
rect 501294 471044 501394 471144
rect 500398 470820 500498 470920
rect 500622 470820 500722 470920
rect 500846 470820 500946 470920
rect 501070 470820 501170 470920
rect 501294 470820 501394 470920
rect 500398 470596 500498 470696
rect 500622 470596 500722 470696
rect 500846 470596 500946 470696
rect 501070 470596 501170 470696
rect 501294 470596 501394 470696
rect 500398 470372 500498 470472
rect 500622 470372 500722 470472
rect 500846 470372 500946 470472
rect 501070 470372 501170 470472
rect 501294 470372 501394 470472
rect 506376 470430 506428 470482
rect 500398 470148 500498 470248
rect 500622 470148 500722 470248
rect 500846 470148 500946 470248
rect 501070 470148 501170 470248
rect 501294 470148 501394 470248
rect 502874 470140 502978 470192
rect 509940 470124 510010 470184
rect 510034 470124 510104 470184
rect 500398 469924 500498 470024
rect 500622 469924 500722 470024
rect 500846 469924 500946 470024
rect 501070 469924 501170 470024
rect 501294 469924 501394 470024
rect 509940 470052 510010 470112
rect 510034 470052 510104 470112
rect 509940 469980 510010 470040
rect 510034 469980 510104 470040
rect 509940 469908 510010 469968
rect 510034 469908 510104 469968
rect 500398 469700 500498 469800
rect 500622 469700 500722 469800
rect 500846 469700 500946 469800
rect 501070 469700 501170 469800
rect 501294 469700 501394 469800
rect 502670 469682 502784 469876
rect 506370 469682 506428 469876
rect 509940 469836 510010 469896
rect 510034 469836 510104 469896
rect 509940 469764 510010 469824
rect 510034 469764 510104 469824
rect 509940 469692 510010 469752
rect 510034 469692 510104 469752
rect 509940 469620 510010 469680
rect 510034 469620 510104 469680
rect 500398 469476 500498 469576
rect 500622 469476 500722 469576
rect 500846 469476 500946 469576
rect 501070 469476 501170 469576
rect 501294 469476 501394 469576
rect 502874 469518 502978 469570
rect 500398 469252 500498 469352
rect 500622 469252 500722 469352
rect 500846 469252 500946 469352
rect 501070 469252 501170 469352
rect 501294 469252 501394 469352
rect 500398 469028 500498 469128
rect 500622 469028 500722 469128
rect 500846 469028 500946 469128
rect 501070 469028 501170 469128
rect 501294 469028 501394 469128
rect 502874 469060 502978 469112
rect 502674 468944 502778 468996
rect 500398 468804 500498 468904
rect 500622 468804 500722 468904
rect 500846 468804 500946 468904
rect 501070 468804 501170 468904
rect 501294 468804 501394 468904
rect 500398 468580 500498 468680
rect 500622 468580 500722 468680
rect 500846 468580 500946 468680
rect 501070 468580 501170 468680
rect 501294 468580 501394 468680
rect 505802 468668 506056 468720
rect 502874 468484 502978 468536
rect 500398 468356 500498 468456
rect 500622 468356 500722 468456
rect 500846 468356 500946 468456
rect 501070 468356 501170 468456
rect 501294 468356 501394 468456
rect 502674 468372 502778 468424
rect 500398 468132 500498 468232
rect 500622 468132 500722 468232
rect 500846 468132 500946 468232
rect 501070 468132 501170 468232
rect 501294 468132 501394 468232
rect 505802 468108 506056 468160
rect 500398 467908 500498 468008
rect 500622 467908 500722 468008
rect 500846 467908 500946 468008
rect 501070 467908 501170 468008
rect 501294 467908 501394 468008
rect 502874 467912 502978 467964
rect 502674 467800 502778 467852
rect 500398 467684 500498 467784
rect 500622 467684 500722 467784
rect 500846 467684 500946 467784
rect 501070 467684 501170 467784
rect 501294 467684 501394 467784
rect 505802 467548 506056 467600
rect 502874 467340 502978 467392
rect 505708 467118 505766 467122
rect 505708 466934 505715 467118
rect 505715 466934 505749 467118
rect 505749 466934 505766 467118
rect 505708 466914 505766 466934
rect 508218 466944 508272 467088
rect 502874 466768 502978 466820
rect 506102 466768 506206 466820
rect 505802 466648 506056 466700
rect 505704 466546 505762 466550
rect 505704 466362 505715 466546
rect 505715 466362 505749 466546
rect 505749 466362 505762 466546
rect 505704 466342 505762 466362
rect 508358 466372 508412 466516
rect 502874 466196 502978 466248
rect 506102 466196 506206 466248
rect 505708 465974 505766 465978
rect 505708 465790 505715 465974
rect 505715 465790 505749 465974
rect 505749 465790 505766 465974
rect 505708 465770 505766 465790
rect 508218 465800 508272 465944
rect 502874 465624 502978 465676
rect 506102 465624 506206 465676
rect 505802 465504 506056 465556
rect 505708 465402 505766 465406
rect 505708 465218 505715 465402
rect 505715 465218 505749 465402
rect 505749 465218 505766 465402
rect 505708 465198 505766 465218
rect 508358 465228 508412 465372
rect 502874 465052 502978 465104
rect 506102 465052 506206 465104
rect 505708 464830 505766 464834
rect 505708 464646 505715 464830
rect 505715 464646 505749 464830
rect 505749 464646 505766 464830
rect 505708 464626 505766 464646
rect 508218 464656 508272 464800
rect 502874 464480 502978 464532
rect 506102 464480 506206 464532
rect 505802 464360 506056 464412
rect 505708 464258 505766 464262
rect 505708 464074 505715 464258
rect 505715 464074 505749 464258
rect 505749 464074 505766 464258
rect 505708 464054 505766 464074
rect 508358 464084 508412 464228
rect 502874 463908 502978 463960
rect 506102 463908 506206 463960
rect 500398 463710 500498 463810
rect 500622 463710 500722 463810
rect 500846 463710 500946 463810
rect 501070 463710 501170 463810
rect 501294 463710 501394 463810
rect 502674 463796 502778 463848
rect 500398 463486 500498 463586
rect 500622 463486 500722 463586
rect 500846 463486 500946 463586
rect 501070 463486 501170 463586
rect 501294 463486 501394 463586
rect 505802 463560 506056 463612
rect 500398 463262 500498 463362
rect 500622 463262 500722 463362
rect 500846 463262 500946 463362
rect 501070 463262 501170 463362
rect 501294 463262 501394 463362
rect 502874 463336 502978 463388
rect 502674 463224 502778 463276
rect 500398 463038 500498 463138
rect 500622 463038 500722 463138
rect 500846 463038 500946 463138
rect 501070 463038 501170 463138
rect 501294 463038 501394 463138
rect 505802 463000 506056 463052
rect 500398 462814 500498 462914
rect 500622 462814 500722 462914
rect 500846 462814 500946 462914
rect 501070 462814 501170 462914
rect 501294 462814 501394 462914
rect 502874 462764 502978 462816
rect 500398 462590 500498 462690
rect 500622 462590 500722 462690
rect 500846 462590 500946 462690
rect 501070 462590 501170 462690
rect 501294 462590 501394 462690
rect 502674 462652 502778 462704
rect 500398 462366 500498 462466
rect 500622 462366 500722 462466
rect 500846 462366 500946 462466
rect 501070 462366 501170 462466
rect 501294 462366 501394 462466
rect 505802 462440 506056 462492
rect 500398 462142 500498 462242
rect 500622 462142 500722 462242
rect 500846 462142 500946 462242
rect 501070 462142 501170 462242
rect 501294 462142 501394 462242
rect 502874 462192 502978 462244
rect 502874 462082 502978 462134
rect 500398 461918 500498 462018
rect 500622 461918 500722 462018
rect 500846 461918 500946 462018
rect 501070 461918 501170 462018
rect 501294 461918 501394 462018
rect 500398 461694 500498 461794
rect 500622 461694 500722 461794
rect 500846 461694 500946 461794
rect 501070 461694 501170 461794
rect 501294 461694 501394 461794
rect 502874 461624 502978 461676
rect 500398 461470 500498 461570
rect 500622 461470 500722 461570
rect 500846 461470 500946 461570
rect 501070 461470 501170 461570
rect 501294 461470 501394 461570
rect 500398 461246 500498 461346
rect 500622 461246 500722 461346
rect 500846 461246 500946 461346
rect 501070 461246 501170 461346
rect 501294 461246 501394 461346
rect 508212 461200 508292 461310
rect 511532 461190 511824 461310
rect 525666 472484 526492 472498
rect 525666 461268 525680 472484
rect 525680 461268 526478 472484
rect 526478 461268 526492 472484
rect 525666 461254 526492 461268
rect 527618 472388 527718 472488
rect 527842 472388 527942 472488
rect 528066 472388 528166 472488
rect 528290 472388 528390 472488
rect 528514 472388 528614 472488
rect 527618 472164 527718 472264
rect 527842 472164 527942 472264
rect 528066 472164 528166 472264
rect 528290 472164 528390 472264
rect 528514 472164 528614 472264
rect 527618 471940 527718 472040
rect 527842 471940 527942 472040
rect 528066 471940 528166 472040
rect 528290 471940 528390 472040
rect 528514 471940 528614 472040
rect 527618 471716 527718 471816
rect 527842 471716 527942 471816
rect 528066 471716 528166 471816
rect 528290 471716 528390 471816
rect 528514 471716 528614 471816
rect 527618 471492 527718 471592
rect 527842 471492 527942 471592
rect 528066 471492 528166 471592
rect 528290 471492 528390 471592
rect 528514 471492 528614 471592
rect 527618 471268 527718 471368
rect 527842 471268 527942 471368
rect 528066 471268 528166 471368
rect 528290 471268 528390 471368
rect 528514 471268 528614 471368
rect 527618 471044 527718 471144
rect 527842 471044 527942 471144
rect 528066 471044 528166 471144
rect 528290 471044 528390 471144
rect 528514 471044 528614 471144
rect 527618 470820 527718 470920
rect 527842 470820 527942 470920
rect 528066 470820 528166 470920
rect 528290 470820 528390 470920
rect 528514 470820 528614 470920
rect 527618 470596 527718 470696
rect 527842 470596 527942 470696
rect 528066 470596 528166 470696
rect 528290 470596 528390 470696
rect 528514 470596 528614 470696
rect 527618 470372 527718 470472
rect 527842 470372 527942 470472
rect 528066 470372 528166 470472
rect 528290 470372 528390 470472
rect 528514 470372 528614 470472
rect 527618 470148 527718 470248
rect 527842 470148 527942 470248
rect 528066 470148 528166 470248
rect 528290 470148 528390 470248
rect 528514 470148 528614 470248
rect 527618 469924 527718 470024
rect 527842 469924 527942 470024
rect 528066 469924 528166 470024
rect 528290 469924 528390 470024
rect 528514 469924 528614 470024
rect 527618 469700 527718 469800
rect 527842 469700 527942 469800
rect 528066 469700 528166 469800
rect 528290 469700 528390 469800
rect 528514 469700 528614 469800
rect 527618 469476 527718 469576
rect 527842 469476 527942 469576
rect 528066 469476 528166 469576
rect 528290 469476 528390 469576
rect 528514 469476 528614 469576
rect 527618 469252 527718 469352
rect 527842 469252 527942 469352
rect 528066 469252 528166 469352
rect 528290 469252 528390 469352
rect 528514 469252 528614 469352
rect 527618 469028 527718 469128
rect 527842 469028 527942 469128
rect 528066 469028 528166 469128
rect 528290 469028 528390 469128
rect 528514 469028 528614 469128
rect 527618 468804 527718 468904
rect 527842 468804 527942 468904
rect 528066 468804 528166 468904
rect 528290 468804 528390 468904
rect 528514 468804 528614 468904
rect 527618 468580 527718 468680
rect 527842 468580 527942 468680
rect 528066 468580 528166 468680
rect 528290 468580 528390 468680
rect 528514 468580 528614 468680
rect 527618 468356 527718 468456
rect 527842 468356 527942 468456
rect 528066 468356 528166 468456
rect 528290 468356 528390 468456
rect 528514 468356 528614 468456
rect 527618 468132 527718 468232
rect 527842 468132 527942 468232
rect 528066 468132 528166 468232
rect 528290 468132 528390 468232
rect 528514 468132 528614 468232
rect 527618 467908 527718 468008
rect 527842 467908 527942 468008
rect 528066 467908 528166 468008
rect 528290 467908 528390 468008
rect 528514 467908 528614 468008
rect 527618 467684 527718 467784
rect 527842 467684 527942 467784
rect 528066 467684 528166 467784
rect 528290 467684 528390 467784
rect 528514 467684 528614 467784
rect 527618 463710 527718 463810
rect 527842 463710 527942 463810
rect 528066 463710 528166 463810
rect 528290 463710 528390 463810
rect 528514 463710 528614 463810
rect 527618 463486 527718 463586
rect 527842 463486 527942 463586
rect 528066 463486 528166 463586
rect 528290 463486 528390 463586
rect 528514 463486 528614 463586
rect 527618 463262 527718 463362
rect 527842 463262 527942 463362
rect 528066 463262 528166 463362
rect 528290 463262 528390 463362
rect 528514 463262 528614 463362
rect 527618 463038 527718 463138
rect 527842 463038 527942 463138
rect 528066 463038 528166 463138
rect 528290 463038 528390 463138
rect 528514 463038 528614 463138
rect 527618 462814 527718 462914
rect 527842 462814 527942 462914
rect 528066 462814 528166 462914
rect 528290 462814 528390 462914
rect 528514 462814 528614 462914
rect 527618 462590 527718 462690
rect 527842 462590 527942 462690
rect 528066 462590 528166 462690
rect 528290 462590 528390 462690
rect 528514 462590 528614 462690
rect 527618 462366 527718 462466
rect 527842 462366 527942 462466
rect 528066 462366 528166 462466
rect 528290 462366 528390 462466
rect 528514 462366 528614 462466
rect 527618 462142 527718 462242
rect 527842 462142 527942 462242
rect 528066 462142 528166 462242
rect 528290 462142 528390 462242
rect 528514 462142 528614 462242
rect 527618 461918 527718 462018
rect 527842 461918 527942 462018
rect 528066 461918 528166 462018
rect 528290 461918 528390 462018
rect 528514 461918 528614 462018
rect 527618 461694 527718 461794
rect 527842 461694 527942 461794
rect 528066 461694 528166 461794
rect 528290 461694 528390 461794
rect 528514 461694 528614 461794
rect 527618 461470 527718 461570
rect 527842 461470 527942 461570
rect 528066 461470 528166 461570
rect 528290 461470 528390 461570
rect 528514 461470 528614 461570
rect 527618 461246 527718 461346
rect 527842 461246 527942 461346
rect 528066 461246 528166 461346
rect 528290 461246 528390 461346
rect 528514 461246 528614 461346
rect 500398 461022 500498 461122
rect 500622 461022 500722 461122
rect 500846 461022 500946 461122
rect 501070 461022 501170 461122
rect 501294 461022 501394 461122
rect 502874 461012 502978 461064
rect 527618 461022 527718 461122
rect 527842 461022 527942 461122
rect 528066 461022 528166 461122
rect 528290 461022 528390 461122
rect 528514 461022 528614 461122
rect 500398 460798 500498 460898
rect 500622 460798 500722 460898
rect 500846 460798 500946 460898
rect 501070 460798 501170 460898
rect 501294 460798 501394 460898
rect 508352 460734 508432 460854
rect 512116 460734 512530 460854
rect 527618 460798 527718 460898
rect 527842 460798 527942 460898
rect 528066 460798 528166 460898
rect 528290 460798 528390 460898
rect 528514 460798 528614 460898
rect 500398 460574 500498 460674
rect 500622 460574 500722 460674
rect 500846 460574 500946 460674
rect 501070 460574 501170 460674
rect 501294 460574 501394 460674
rect 527618 460574 527718 460674
rect 527842 460574 527942 460674
rect 528066 460574 528166 460674
rect 528290 460574 528390 460674
rect 528514 460574 528614 460674
rect 500398 460350 500498 460450
rect 500622 460350 500722 460450
rect 500846 460350 500946 460450
rect 501070 460350 501170 460450
rect 501294 460350 501394 460450
rect 500398 460126 500498 460226
rect 500622 460126 500722 460226
rect 500846 460126 500946 460226
rect 501070 460126 501170 460226
rect 501294 460126 501394 460226
rect 500398 459902 500498 460002
rect 500622 459902 500722 460002
rect 500846 459902 500946 460002
rect 501070 459902 501170 460002
rect 501294 459902 501394 460002
rect 500398 459678 500498 459778
rect 500622 459678 500722 459778
rect 500846 459678 500946 459778
rect 501070 459678 501170 459778
rect 501294 459678 501394 459778
rect 500398 459454 500498 459554
rect 500622 459454 500722 459554
rect 500846 459454 500946 459554
rect 501070 459454 501170 459554
rect 501294 459454 501394 459554
rect 500398 459230 500498 459330
rect 500622 459230 500722 459330
rect 500846 459230 500946 459330
rect 501070 459230 501170 459330
rect 501294 459230 501394 459330
rect 502528 459952 502628 460352
rect 502814 459974 502962 460442
rect 505802 459974 506056 460442
rect 527618 460350 527718 460450
rect 527842 460350 527942 460450
rect 528066 460350 528166 460450
rect 528290 460350 528390 460450
rect 528514 460350 528614 460450
rect 527618 460126 527718 460226
rect 527842 460126 527942 460226
rect 528066 460126 528166 460226
rect 528290 460126 528390 460226
rect 528514 460126 528614 460226
rect 527618 459902 527718 460002
rect 527842 459902 527942 460002
rect 528066 459902 528166 460002
rect 528290 459902 528390 460002
rect 528514 459902 528614 460002
rect 500398 459006 500498 459106
rect 500622 459006 500722 459106
rect 500846 459006 500946 459106
rect 501070 459006 501170 459106
rect 501294 459006 501394 459106
rect 502828 458982 502948 459122
rect 500398 458782 500498 458882
rect 500622 458782 500722 458882
rect 500846 458782 500946 458882
rect 501070 458782 501170 458882
rect 501294 458782 501394 458882
rect 502668 458782 502748 458862
rect 500398 458558 500498 458658
rect 500622 458558 500722 458658
rect 500846 458558 500946 458658
rect 501070 458558 501170 458658
rect 501294 458558 501394 458658
rect 502828 458522 502948 458662
rect 500398 458334 500498 458434
rect 500622 458334 500722 458434
rect 500846 458334 500946 458434
rect 501070 458334 501170 458434
rect 501294 458334 501394 458434
rect 500398 458110 500498 458210
rect 500622 458110 500722 458210
rect 500846 458110 500946 458210
rect 501070 458110 501170 458210
rect 501294 458110 501394 458210
rect 502828 458062 502948 458202
rect 500398 457886 500498 457986
rect 500622 457886 500722 457986
rect 500846 457886 500946 457986
rect 501070 457886 501170 457986
rect 501294 457886 501394 457986
rect 502668 457862 502748 457942
rect 500398 457662 500498 457762
rect 500622 457662 500722 457762
rect 500846 457662 500946 457762
rect 501070 457662 501170 457762
rect 501294 457662 501394 457762
rect 502828 457602 502948 457742
rect 500398 457438 500498 457538
rect 500622 457438 500722 457538
rect 500846 457438 500946 457538
rect 501070 457438 501170 457538
rect 501294 457438 501394 457538
rect 512134 457348 512422 459336
rect 512836 457348 513286 459336
rect 527618 459678 527718 459778
rect 527842 459678 527942 459778
rect 528066 459678 528166 459778
rect 528290 459678 528390 459778
rect 528514 459678 528614 459778
rect 527618 459454 527718 459554
rect 527842 459454 527942 459554
rect 528066 459454 528166 459554
rect 528290 459454 528390 459554
rect 528514 459454 528614 459554
rect 527618 459230 527718 459330
rect 527842 459230 527942 459330
rect 528066 459230 528166 459330
rect 528290 459230 528390 459330
rect 528514 459230 528614 459330
rect 527618 459006 527718 459106
rect 527842 459006 527942 459106
rect 528066 459006 528166 459106
rect 528290 459006 528390 459106
rect 528514 459006 528614 459106
rect 527618 458782 527718 458882
rect 527842 458782 527942 458882
rect 528066 458782 528166 458882
rect 528290 458782 528390 458882
rect 528514 458782 528614 458882
rect 527618 458558 527718 458658
rect 527842 458558 527942 458658
rect 528066 458558 528166 458658
rect 528290 458558 528390 458658
rect 528514 458558 528614 458658
rect 500398 457214 500498 457314
rect 500622 457214 500722 457314
rect 500846 457214 500946 457314
rect 501070 457214 501170 457314
rect 501294 457214 501394 457314
rect 502828 457142 502948 457282
rect 502668 456942 502748 457022
rect 502828 456682 502948 456822
rect 502828 456222 502948 456362
rect 502668 456022 502748 456102
rect 502828 455762 502948 455902
rect 502828 455302 502948 455442
rect 502668 455102 502748 455182
rect 502828 454842 502948 454982
rect 511534 454648 511822 456636
rect 502528 454042 502628 454442
rect 502828 453482 502948 453622
rect 513720 453556 513920 453756
rect 514154 453556 514354 453756
rect 514588 453556 514788 453756
rect 502668 453282 502748 453362
rect 502828 453022 502948 453162
rect 513720 453122 513920 453322
rect 514154 453122 514354 453322
rect 514588 453122 514788 453322
rect 502828 452562 502948 452702
rect 513720 452688 513920 452888
rect 514154 452688 514354 452888
rect 514588 452688 514788 452888
rect 502668 452362 502748 452442
rect 502828 452102 502948 452242
rect 513720 452254 513920 452454
rect 514154 452254 514354 452454
rect 514588 452254 514788 452454
rect 513720 451820 513920 452020
rect 514154 451820 514354 452020
rect 514588 451820 514788 452020
rect 502828 451642 502948 451782
rect 502668 451442 502748 451522
rect 513720 451386 513920 451586
rect 514154 451386 514354 451586
rect 514588 451386 514788 451586
rect 502828 451182 502948 451322
rect 513720 450952 513920 451152
rect 514154 450952 514354 451152
rect 514588 450952 514788 451152
rect 502828 450722 502948 450862
rect 502668 450522 502748 450602
rect 513720 450518 513920 450718
rect 514154 450518 514354 450718
rect 514588 450518 514788 450718
rect 502828 450262 502948 450402
rect 513720 450084 513920 450284
rect 514154 450084 514354 450284
rect 514588 450084 514788 450284
rect 502828 449802 502948 449942
rect 502668 449602 502748 449682
rect 513720 449650 513920 449850
rect 514154 449650 514354 449850
rect 514588 449650 514788 449850
rect 502828 449342 502948 449482
rect 513720 449216 513920 449416
rect 514154 449216 514354 449416
rect 514588 449216 514788 449416
rect 502528 448542 502628 448942
rect 514588 448816 514788 449016
rect 514588 448416 514788 448616
rect 502828 447982 502948 448122
rect 502668 447782 502748 447862
rect 502828 447522 502948 447662
rect 502828 447062 502948 447202
rect 502668 446862 502748 446942
rect 502828 446602 502948 446742
rect 511534 446348 511822 448336
rect 514588 448016 514788 448216
rect 515396 450322 515954 450880
rect 516196 450870 516616 450880
rect 516196 450332 516207 450870
rect 516207 450332 516605 450870
rect 516605 450332 516616 450870
rect 516196 450322 516616 450332
rect 516196 450052 516616 450062
rect 516196 449514 516208 450052
rect 516208 449514 516605 450052
rect 516605 449514 516616 450052
rect 516196 449504 516616 449514
rect 516196 449234 516616 449244
rect 516196 448696 516208 449234
rect 516208 448696 516605 449234
rect 516605 448696 516616 449234
rect 516196 448686 516616 448696
rect 527618 458334 527718 458434
rect 527842 458334 527942 458434
rect 528066 458334 528166 458434
rect 528290 458334 528390 458434
rect 528514 458334 528614 458434
rect 527618 458110 527718 458210
rect 527842 458110 527942 458210
rect 528066 458110 528166 458210
rect 528290 458110 528390 458210
rect 528514 458110 528614 458210
rect 527618 457886 527718 457986
rect 527842 457886 527942 457986
rect 528066 457886 528166 457986
rect 528290 457886 528390 457986
rect 528514 457886 528614 457986
rect 527618 457662 527718 457762
rect 527842 457662 527942 457762
rect 528066 457662 528166 457762
rect 528290 457662 528390 457762
rect 528514 457662 528614 457762
rect 527618 457438 527718 457538
rect 527842 457438 527942 457538
rect 528066 457438 528166 457538
rect 528290 457438 528390 457538
rect 528514 457438 528614 457538
rect 527618 457214 527718 457314
rect 527842 457214 527942 457314
rect 528066 457214 528166 457314
rect 528290 457214 528390 457314
rect 528514 457214 528614 457314
rect 522994 455778 523414 455788
rect 522994 455240 523005 455778
rect 523005 455240 523402 455778
rect 523402 455240 523414 455778
rect 522994 455230 523414 455240
rect 523594 455230 524152 455788
rect 522198 454412 522690 454970
rect 522994 454960 523414 454970
rect 522994 454422 523005 454960
rect 523005 454422 523402 454960
rect 523402 454422 523414 454960
rect 522994 454412 523414 454422
rect 522132 450322 522690 450880
rect 522932 450870 523352 450880
rect 522932 450332 522943 450870
rect 522943 450332 523340 450870
rect 523340 450332 523352 450870
rect 522932 450322 523352 450332
rect 516858 448686 517416 449244
rect 517658 449504 518216 450062
rect 515396 447868 515954 448426
rect 516196 448416 516616 448426
rect 516196 447878 516207 448416
rect 516207 447878 516605 448416
rect 516605 447878 516616 448416
rect 516196 447868 516616 447878
rect 514588 447616 514788 447816
rect 514588 447216 514788 447416
rect 516196 447598 516616 447608
rect 516196 447060 516208 447598
rect 516208 447060 516605 447598
rect 516605 447060 516616 447598
rect 516196 447050 516616 447060
rect 516858 447050 517416 447608
rect 514588 446816 514788 447016
rect 514588 446416 514788 446616
rect 502828 446142 502948 446282
rect 516196 446780 516616 446790
rect 516196 446242 516208 446780
rect 516208 446242 516605 446780
rect 516605 446242 516616 446780
rect 516196 446232 516616 446242
rect 502668 445942 502748 446022
rect 514588 446016 514788 446216
rect 502828 445682 502948 445822
rect 502828 445222 502948 445362
rect 502668 445022 502748 445102
rect 502828 444762 502948 444902
rect 502828 444302 502948 444442
rect 502668 444102 502748 444182
rect 502828 443842 502948 443982
rect 512134 443648 512422 445636
rect 512836 443648 513286 445636
rect 514588 445616 514788 445816
rect 514588 444016 514788 444216
rect 514588 443616 514788 443816
rect 514588 443216 514788 443416
rect 502526 442586 502626 442986
rect 514588 442816 514788 443016
rect 514588 442416 514788 442616
rect 514588 442016 514788 442216
rect 515396 445414 515954 445972
rect 516196 445962 516616 445972
rect 516196 445424 516207 445962
rect 516207 445424 516605 445962
rect 516605 445424 516616 445962
rect 516196 445414 516616 445424
rect 516066 445154 516584 445232
rect 516066 445144 516616 445154
rect 516066 444606 516208 445144
rect 516208 444606 516605 445144
rect 516605 444606 516616 445144
rect 516066 444596 516616 444606
rect 516066 444540 516584 444596
rect 516196 444326 516616 444336
rect 516196 443788 516208 444326
rect 516208 443788 516605 444326
rect 516605 443788 516616 444326
rect 516196 443778 516616 443788
rect 516196 443508 516616 443518
rect 516196 442970 516208 443508
rect 516208 442970 516605 443508
rect 516605 442970 516616 443508
rect 516196 442960 516616 442970
rect 522932 450052 523352 450062
rect 522932 449514 522943 450052
rect 522943 449514 523340 450052
rect 523340 449514 523352 450052
rect 522932 449504 523352 449514
rect 562480 455360 562560 455440
rect 562640 455360 562720 455440
rect 562800 455360 562880 455440
rect 562960 455360 563040 455440
rect 563120 455360 563200 455440
rect 563280 455360 563360 455440
rect 563440 455360 563520 455440
rect 563600 455360 563680 455440
rect 563760 455360 563840 455440
rect 563920 455360 564000 455440
rect 564080 455360 564160 455440
rect 564240 455360 564320 455440
rect 564400 455360 564480 455440
rect 564560 455360 564640 455440
rect 564720 455360 564800 455440
rect 564880 455360 564960 455440
rect 565040 455360 565120 455440
rect 565200 455360 565280 455440
rect 565360 455360 565440 455440
rect 565520 455360 565600 455440
rect 565680 455360 565760 455440
rect 565840 455360 565920 455440
rect 566000 455360 566080 455440
rect 566160 455360 566240 455440
rect 566320 455360 566400 455440
rect 566480 455360 566560 455440
rect 566640 455360 566720 455440
rect 566800 455360 566880 455440
rect 566960 455360 567040 455440
rect 567120 455360 567200 455440
rect 567280 455360 567360 455440
rect 562480 455212 562560 455280
rect 562640 455212 562720 455280
rect 562800 455212 562880 455280
rect 562960 455212 563040 455280
rect 563120 455212 563200 455280
rect 563280 455212 563360 455280
rect 563440 455212 563520 455280
rect 563600 455212 563680 455280
rect 563760 455212 563840 455280
rect 563920 455212 564000 455280
rect 564080 455212 564160 455280
rect 564240 455212 564320 455280
rect 564400 455212 564480 455280
rect 564560 455212 564640 455280
rect 564720 455212 564800 455280
rect 564880 455212 564960 455280
rect 565040 455212 565120 455280
rect 565200 455212 565280 455280
rect 565360 455212 565440 455280
rect 565520 455212 565600 455280
rect 565680 455212 565760 455280
rect 565840 455212 565920 455280
rect 566000 455212 566080 455280
rect 566160 455212 566240 455280
rect 566320 455212 566400 455280
rect 566480 455212 566560 455280
rect 566640 455212 566720 455280
rect 566800 455212 566880 455280
rect 566960 455212 567040 455280
rect 567120 455212 567200 455280
rect 567280 455212 567360 455280
rect 562480 455200 562560 455212
rect 562640 455200 562720 455212
rect 562800 455200 562880 455212
rect 562960 455200 563040 455212
rect 563120 455200 563200 455212
rect 563280 455200 563360 455212
rect 563440 455200 563520 455212
rect 563600 455200 563680 455212
rect 563760 455200 563840 455212
rect 563920 455200 564000 455212
rect 564080 455200 564160 455212
rect 564240 455200 564320 455212
rect 564400 455200 564480 455212
rect 564560 455200 564640 455212
rect 564720 455200 564800 455212
rect 564880 455200 564960 455212
rect 565040 455200 565120 455212
rect 565200 455200 565280 455212
rect 565360 455200 565440 455212
rect 565520 455200 565600 455212
rect 565680 455200 565760 455212
rect 565840 455200 565920 455212
rect 566000 455200 566080 455212
rect 566160 455200 566240 455212
rect 566320 455200 566400 455212
rect 566480 455200 566560 455212
rect 566640 455200 566720 455212
rect 566800 455200 566880 455212
rect 566960 455200 567040 455212
rect 567120 455200 567200 455212
rect 567280 455200 567360 455212
rect 572640 455360 572720 455440
rect 572800 455360 572880 455440
rect 572960 455360 573040 455440
rect 573120 455360 573200 455440
rect 573280 455360 573360 455440
rect 573440 455360 573520 455440
rect 573600 455360 573680 455440
rect 573760 455360 573840 455440
rect 573920 455360 574000 455440
rect 574080 455360 574160 455440
rect 574240 455360 574320 455440
rect 574400 455360 574480 455440
rect 574560 455360 574640 455440
rect 574720 455360 574800 455440
rect 574880 455360 574960 455440
rect 575040 455360 575120 455440
rect 575200 455360 575280 455440
rect 575360 455360 575440 455440
rect 575520 455360 575600 455440
rect 575680 455360 575760 455440
rect 575840 455360 575920 455440
rect 576000 455360 576080 455440
rect 576160 455360 576240 455440
rect 576320 455360 576400 455440
rect 576480 455360 576560 455440
rect 576640 455360 576720 455440
rect 576800 455360 576880 455440
rect 576960 455360 577040 455440
rect 577120 455360 577200 455440
rect 577280 455360 577360 455440
rect 577440 455360 577520 455440
rect 572640 455246 572720 455280
rect 572800 455246 572880 455280
rect 572960 455246 573040 455280
rect 573120 455246 573200 455280
rect 573280 455246 573360 455280
rect 573440 455246 573520 455280
rect 573600 455246 573680 455280
rect 573760 455246 573840 455280
rect 573920 455246 574000 455280
rect 574080 455246 574160 455280
rect 574240 455246 574320 455280
rect 574400 455246 574480 455280
rect 574560 455246 574640 455280
rect 574720 455246 574800 455280
rect 574880 455246 574960 455280
rect 575040 455246 575120 455280
rect 575200 455246 575280 455280
rect 575360 455246 575440 455280
rect 575520 455246 575600 455280
rect 575680 455246 575760 455280
rect 575840 455246 575920 455280
rect 576000 455246 576080 455280
rect 576160 455246 576240 455280
rect 576320 455246 576400 455280
rect 576480 455246 576560 455280
rect 576640 455246 576720 455280
rect 576800 455246 576880 455280
rect 576960 455246 577040 455280
rect 577120 455246 577200 455280
rect 577280 455246 577360 455280
rect 577440 455246 577520 455280
rect 572640 455212 572720 455246
rect 572800 455212 572880 455246
rect 572960 455212 573040 455246
rect 573120 455212 573200 455246
rect 573280 455212 573360 455246
rect 573440 455212 573520 455246
rect 573600 455212 573680 455246
rect 573760 455212 573840 455246
rect 573920 455212 574000 455246
rect 574080 455212 574160 455246
rect 574240 455212 574320 455246
rect 574400 455212 574480 455246
rect 574560 455212 574640 455246
rect 574720 455212 574800 455246
rect 574880 455212 574960 455246
rect 575040 455212 575120 455246
rect 575200 455212 575280 455246
rect 575360 455212 575440 455246
rect 575520 455212 575600 455246
rect 575680 455212 575760 455246
rect 575840 455212 575920 455246
rect 576000 455212 576080 455246
rect 576160 455212 576240 455246
rect 576320 455212 576400 455246
rect 576480 455212 576560 455246
rect 576640 455212 576720 455246
rect 576800 455212 576880 455246
rect 576960 455212 577040 455246
rect 577120 455212 577200 455246
rect 577280 455212 577360 455246
rect 577440 455212 577520 455246
rect 572640 455200 572720 455212
rect 572800 455200 572880 455212
rect 572960 455200 573040 455212
rect 573120 455200 573200 455212
rect 573280 455200 573360 455212
rect 573440 455200 573520 455212
rect 573600 455200 573680 455212
rect 573760 455200 573840 455212
rect 573920 455200 574000 455212
rect 574080 455200 574160 455212
rect 574240 455200 574320 455212
rect 574400 455200 574480 455212
rect 574560 455200 574640 455212
rect 574720 455200 574800 455212
rect 574880 455200 574960 455212
rect 575040 455200 575120 455212
rect 575200 455200 575280 455212
rect 575360 455200 575440 455212
rect 575520 455200 575600 455212
rect 575680 455200 575760 455212
rect 575840 455200 575920 455212
rect 576000 455200 576080 455212
rect 576160 455200 576240 455212
rect 576320 455200 576400 455212
rect 576480 455200 576560 455212
rect 576640 455200 576720 455212
rect 576800 455200 576880 455212
rect 576960 455200 577040 455212
rect 577120 455200 577200 455212
rect 577280 455200 577360 455212
rect 577440 455200 577520 455212
rect 562222 453859 562282 453919
rect 562342 453859 562402 453919
rect 562462 453859 562522 453919
rect 562582 453859 562642 453919
rect 562702 453859 562762 453919
rect 562822 453859 562882 453919
rect 562942 453859 563002 453919
rect 563062 453859 563122 453919
rect 563182 453859 563242 453919
rect 563302 453859 563362 453919
rect 563422 453859 563482 453919
rect 563542 453859 563602 453919
rect 563662 453859 563722 453919
rect 563782 453859 563842 453919
rect 563902 453859 563962 453919
rect 564022 453859 564082 453919
rect 564142 453859 564202 453919
rect 564262 453859 564322 453919
rect 564382 453859 564442 453919
rect 564502 453859 564562 453919
rect 564622 453859 564682 453919
rect 564742 453859 564802 453919
rect 564862 453859 564922 453919
rect 564982 453859 565042 453919
rect 565102 453859 565162 453919
rect 565222 453859 565282 453919
rect 565342 453859 565402 453919
rect 565462 453859 565522 453919
rect 565582 453859 565642 453919
rect 565702 453859 565762 453919
rect 565822 453859 565882 453919
rect 565942 453859 566002 453919
rect 566062 453859 566122 453919
rect 566182 453859 566242 453919
rect 566302 453859 566362 453919
rect 566422 453859 566482 453919
rect 566542 453859 566602 453919
rect 566662 453859 566722 453919
rect 566782 453859 566842 453919
rect 566902 453859 566962 453919
rect 567022 453859 567082 453919
rect 567142 453859 567202 453919
rect 567262 453859 567322 453919
rect 567382 453859 567442 453919
rect 567502 453859 567562 453919
rect 562222 453739 562282 453799
rect 562342 453739 562402 453799
rect 562462 453739 562522 453799
rect 562582 453739 562642 453799
rect 562702 453739 562762 453799
rect 562822 453739 562882 453799
rect 562942 453739 563002 453799
rect 563062 453739 563122 453799
rect 563182 453739 563242 453799
rect 563302 453739 563362 453799
rect 563422 453739 563482 453799
rect 563542 453739 563602 453799
rect 563662 453739 563722 453799
rect 563782 453739 563842 453799
rect 563902 453739 563962 453799
rect 564022 453739 564082 453799
rect 564142 453739 564202 453799
rect 564262 453739 564322 453799
rect 564382 453739 564442 453799
rect 564502 453739 564562 453799
rect 564622 453739 564682 453799
rect 564742 453739 564802 453799
rect 564862 453739 564922 453799
rect 564982 453739 565042 453799
rect 565102 453739 565162 453799
rect 565222 453739 565282 453799
rect 565342 453739 565402 453799
rect 565462 453739 565522 453799
rect 565582 453739 565642 453799
rect 565702 453739 565762 453799
rect 565822 453739 565882 453799
rect 565942 453739 566002 453799
rect 566062 453739 566122 453799
rect 566182 453739 566242 453799
rect 566302 453739 566362 453799
rect 566422 453739 566482 453799
rect 566542 453739 566602 453799
rect 566662 453739 566722 453799
rect 566782 453739 566842 453799
rect 566902 453739 566962 453799
rect 567022 453739 567082 453799
rect 567142 453739 567202 453799
rect 567262 453739 567322 453799
rect 567382 453739 567442 453799
rect 567502 453739 567562 453799
rect 572332 453874 572392 453934
rect 572452 453874 572512 453934
rect 572572 453874 572632 453934
rect 572692 453874 572752 453934
rect 572812 453874 572872 453934
rect 572932 453874 572992 453934
rect 573052 453874 573112 453934
rect 573172 453874 573232 453934
rect 573292 453874 573352 453934
rect 573412 453874 573472 453934
rect 573532 453874 573592 453934
rect 573652 453874 573712 453934
rect 573772 453874 573832 453934
rect 573892 453874 573952 453934
rect 574012 453874 574072 453934
rect 574132 453874 574192 453934
rect 574252 453874 574312 453934
rect 574372 453874 574432 453934
rect 574492 453874 574552 453934
rect 574612 453874 574672 453934
rect 574732 453874 574792 453934
rect 574852 453874 574912 453934
rect 574972 453874 575032 453934
rect 575092 453874 575152 453934
rect 575212 453874 575272 453934
rect 575332 453874 575392 453934
rect 575452 453874 575512 453934
rect 575572 453874 575632 453934
rect 575692 453874 575752 453934
rect 575812 453874 575872 453934
rect 575932 453874 575992 453934
rect 576052 453874 576112 453934
rect 576172 453874 576232 453934
rect 576292 453874 576352 453934
rect 576412 453874 576472 453934
rect 576532 453874 576592 453934
rect 576652 453874 576712 453934
rect 576772 453874 576832 453934
rect 576892 453874 576952 453934
rect 577012 453874 577072 453934
rect 577132 453874 577192 453934
rect 577252 453874 577312 453934
rect 577372 453874 577432 453934
rect 577492 453874 577552 453934
rect 577612 453874 577672 453934
rect 572332 453754 572392 453814
rect 572452 453754 572512 453814
rect 572572 453754 572632 453814
rect 572692 453754 572752 453814
rect 572812 453754 572872 453814
rect 572932 453754 572992 453814
rect 573052 453754 573112 453814
rect 573172 453754 573232 453814
rect 573292 453754 573352 453814
rect 573412 453754 573472 453814
rect 573532 453754 573592 453814
rect 573652 453754 573712 453814
rect 573772 453754 573832 453814
rect 573892 453754 573952 453814
rect 574012 453754 574072 453814
rect 574132 453754 574192 453814
rect 574252 453754 574312 453814
rect 574372 453754 574432 453814
rect 574492 453754 574552 453814
rect 574612 453754 574672 453814
rect 574732 453754 574792 453814
rect 574852 453754 574912 453814
rect 574972 453754 575032 453814
rect 575092 453754 575152 453814
rect 575212 453754 575272 453814
rect 575332 453754 575392 453814
rect 575452 453754 575512 453814
rect 575572 453754 575632 453814
rect 575692 453754 575752 453814
rect 575812 453754 575872 453814
rect 575932 453754 575992 453814
rect 576052 453754 576112 453814
rect 576172 453754 576232 453814
rect 576292 453754 576352 453814
rect 576412 453754 576472 453814
rect 576532 453754 576592 453814
rect 576652 453754 576712 453814
rect 576772 453754 576832 453814
rect 576892 453754 576952 453814
rect 577012 453754 577072 453814
rect 577132 453754 577192 453814
rect 577252 453754 577312 453814
rect 577372 453754 577432 453814
rect 577492 453754 577552 453814
rect 577612 453754 577672 453814
rect 523594 449504 524152 450062
rect 522932 449234 523352 449244
rect 522932 448696 522943 449234
rect 522943 448696 523340 449234
rect 523340 448696 523352 449234
rect 522932 448686 523352 448696
rect 524394 448674 524952 449232
rect 517658 446232 518216 446790
rect 522132 447868 522690 448426
rect 522932 448416 523352 448426
rect 522932 447878 522943 448416
rect 522943 447878 523340 448416
rect 523340 447878 523352 448416
rect 522932 447868 523352 447878
rect 522932 447598 523352 447608
rect 522932 447060 522943 447598
rect 522943 447060 523340 447598
rect 523340 447060 523352 447598
rect 522932 447050 523352 447060
rect 524394 447050 524952 447608
rect 522932 446780 523352 446790
rect 522932 446242 522943 446780
rect 522943 446242 523340 446780
rect 523340 446242 523352 446780
rect 522932 446232 523352 446242
rect 523594 446232 524152 446790
rect 522132 445414 522690 445972
rect 522932 445962 523352 445972
rect 522932 445424 522943 445962
rect 522943 445424 523340 445962
rect 523340 445424 523352 445962
rect 522932 445414 523352 445424
rect 522932 445144 523352 445154
rect 522932 444606 522943 445144
rect 522943 444606 523340 445144
rect 523340 444606 523352 445144
rect 522932 444596 523352 444606
rect 516858 442960 517416 443518
rect 517658 443778 518216 444336
rect 515396 442142 515954 442700
rect 516196 442690 516616 442700
rect 516196 442152 516207 442690
rect 516207 442152 516605 442690
rect 516605 442152 516616 442690
rect 516196 442142 516616 442152
rect 503652 440732 504588 441668
rect 513548 440732 514066 441666
rect 514588 441616 514788 441816
rect 514588 441216 514788 441416
rect 516196 441872 516616 441882
rect 516196 441334 516208 441872
rect 516208 441334 516605 441872
rect 516605 441334 516616 441872
rect 516196 441324 516616 441334
rect 522932 444326 523352 444336
rect 522932 443788 522943 444326
rect 522943 443788 523340 444326
rect 523340 443788 523352 444326
rect 522932 443778 523352 443788
rect 523594 443778 524152 444336
rect 522932 443508 523352 443518
rect 522932 442970 522943 443508
rect 522943 442970 523340 443508
rect 523340 442970 523352 443508
rect 522932 442960 523352 442970
rect 524394 442960 524952 443518
rect 517658 441324 518216 441882
rect 522132 442142 522690 442700
rect 515924 441054 516616 441142
rect 514588 440816 514788 441016
rect 515924 440516 516208 441054
rect 516208 440516 516605 441054
rect 516605 440516 516616 441054
rect 515924 440450 516616 440516
rect 508806 439632 509498 440324
rect 512836 439632 513286 440324
rect 515924 440236 516616 440324
rect 515924 439698 516208 440236
rect 516208 439698 516605 440236
rect 516605 439698 516616 440236
rect 515924 439632 516616 439698
rect 522932 442690 523352 442700
rect 522932 442152 522943 442690
rect 522943 442152 523340 442690
rect 523340 442152 523352 442690
rect 522932 442142 523352 442152
rect 522932 441872 523352 441882
rect 522932 441334 522943 441872
rect 522943 441334 523340 441872
rect 523340 441334 523352 441872
rect 522932 441324 523352 441334
rect 523594 441324 524152 441882
rect 522932 441054 523352 441064
rect 522932 440516 522943 441054
rect 522943 440516 523340 441054
rect 523340 440516 523352 441054
rect 522932 440506 523352 440516
rect 522132 439688 522690 440246
rect 522932 440236 523352 440246
rect 522932 439698 522943 440236
rect 522943 439698 523340 440236
rect 523340 439698 523352 440236
rect 522932 439688 523352 439698
rect 511534 438814 511822 439504
rect 515924 439418 516616 439506
rect 515924 438880 516208 439418
rect 516208 438880 516605 439418
rect 516605 438880 516616 439418
rect 515924 438814 516616 438880
rect 522932 439418 523352 439428
rect 522932 438880 522943 439418
rect 522943 438880 523340 439418
rect 523340 438880 523352 439418
rect 522932 438870 523352 438880
rect 524394 440506 524952 441064
rect 523594 438870 524152 439428
rect 500418 437440 500518 437540
rect 500642 437440 500742 437540
rect 500866 437440 500966 437540
rect 501090 437440 501190 437540
rect 501314 437440 501414 437540
rect 500418 437216 500518 437316
rect 500642 437216 500742 437316
rect 500866 437216 500966 437316
rect 501090 437216 501190 437316
rect 501314 437216 501414 437316
rect 500418 436992 500518 437092
rect 500642 436992 500742 437092
rect 500866 436992 500966 437092
rect 501090 436992 501190 437092
rect 501314 436992 501414 437092
rect 500418 436768 500518 436868
rect 500642 436768 500742 436868
rect 500866 436768 500966 436868
rect 501090 436768 501190 436868
rect 501314 436768 501414 436868
rect 500418 436544 500518 436644
rect 500642 436544 500742 436644
rect 500866 436544 500966 436644
rect 501090 436544 501190 436644
rect 501314 436544 501414 436644
rect 500418 436320 500518 436420
rect 500642 436320 500742 436420
rect 500866 436320 500966 436420
rect 501090 436320 501190 436420
rect 501314 436320 501414 436420
rect 500418 436096 500518 436196
rect 500642 436096 500742 436196
rect 500866 436096 500966 436196
rect 501090 436096 501190 436196
rect 501314 436096 501414 436196
rect 500418 435872 500518 435972
rect 500642 435872 500742 435972
rect 500866 435872 500966 435972
rect 501090 435872 501190 435972
rect 501314 435872 501414 435972
rect 500418 435648 500518 435748
rect 500642 435648 500742 435748
rect 500866 435648 500966 435748
rect 501090 435648 501190 435748
rect 501314 435648 501414 435748
rect 500418 435424 500518 435524
rect 500642 435424 500742 435524
rect 500866 435424 500966 435524
rect 501090 435424 501190 435524
rect 501314 435424 501414 435524
rect 500418 435200 500518 435300
rect 500642 435200 500742 435300
rect 500866 435200 500966 435300
rect 501090 435200 501190 435300
rect 501314 435200 501414 435300
rect 500418 434976 500518 435076
rect 500642 434976 500742 435076
rect 500866 434976 500966 435076
rect 501090 434976 501190 435076
rect 501314 434976 501414 435076
rect 500418 434752 500518 434852
rect 500642 434752 500742 434852
rect 500866 434752 500966 434852
rect 501090 434752 501190 434852
rect 501314 434752 501414 434852
rect 500418 434528 500518 434628
rect 500642 434528 500742 434628
rect 500866 434528 500966 434628
rect 501090 434528 501190 434628
rect 501314 434528 501414 434628
rect 500418 434304 500518 434404
rect 500642 434304 500742 434404
rect 500866 434304 500966 434404
rect 501090 434304 501190 434404
rect 501314 434304 501414 434404
rect 500418 434080 500518 434180
rect 500642 434080 500742 434180
rect 500866 434080 500966 434180
rect 501090 434080 501190 434180
rect 501314 434080 501414 434180
rect 500418 433856 500518 433956
rect 500642 433856 500742 433956
rect 500866 433856 500966 433956
rect 501090 433856 501190 433956
rect 501314 433856 501414 433956
rect 500418 433632 500518 433732
rect 500642 433632 500742 433732
rect 500866 433632 500966 433732
rect 501090 433632 501190 433732
rect 501314 433632 501414 433732
rect 500418 433408 500518 433508
rect 500642 433408 500742 433508
rect 500866 433408 500966 433508
rect 501090 433408 501190 433508
rect 501314 433408 501414 433508
rect 500418 433184 500518 433284
rect 500642 433184 500742 433284
rect 500866 433184 500966 433284
rect 501090 433184 501190 433284
rect 501314 433184 501414 433284
rect 500418 432960 500518 433060
rect 500642 432960 500742 433060
rect 500866 432960 500966 433060
rect 501090 432960 501190 433060
rect 501314 432960 501414 433060
rect 500418 432736 500518 432836
rect 500642 432736 500742 432836
rect 500866 432736 500966 432836
rect 501090 432736 501190 432836
rect 501314 432736 501414 432836
rect 500418 432512 500518 432612
rect 500642 432512 500742 432612
rect 500866 432512 500966 432612
rect 501090 432512 501190 432612
rect 501314 432512 501414 432612
rect 500418 432288 500518 432388
rect 500642 432288 500742 432388
rect 500866 432288 500966 432388
rect 501090 432288 501190 432388
rect 501314 432288 501414 432388
rect 503716 436824 503768 436848
rect 503820 436824 503872 436848
rect 503924 436824 503976 436848
rect 503716 436796 503740 436824
rect 503740 436796 503768 436824
rect 503820 436796 503840 436824
rect 503840 436796 503872 436824
rect 503924 436796 503940 436824
rect 503940 436796 503974 436824
rect 503974 436796 503976 436824
rect 504028 436824 504080 436848
rect 504028 436796 504040 436824
rect 504040 436796 504074 436824
rect 504074 436796 504080 436824
rect 504132 436824 504184 436848
rect 504132 436796 504140 436824
rect 504140 436796 504174 436824
rect 504174 436796 504184 436824
rect 504236 436824 504288 436848
rect 504236 436796 504240 436824
rect 504240 436796 504274 436824
rect 504274 436796 504288 436824
rect 503716 436724 503768 436744
rect 503820 436724 503872 436744
rect 503924 436724 503976 436744
rect 503716 436692 503740 436724
rect 503740 436692 503768 436724
rect 503820 436692 503840 436724
rect 503840 436692 503872 436724
rect 503924 436692 503940 436724
rect 503940 436692 503974 436724
rect 503974 436692 503976 436724
rect 504028 436724 504080 436744
rect 504028 436692 504040 436724
rect 504040 436692 504074 436724
rect 504074 436692 504080 436724
rect 504132 436724 504184 436744
rect 504132 436692 504140 436724
rect 504140 436692 504174 436724
rect 504174 436692 504184 436724
rect 504236 436724 504288 436744
rect 504236 436692 504240 436724
rect 504240 436692 504274 436724
rect 504274 436692 504288 436724
rect 503716 436624 503768 436640
rect 503820 436624 503872 436640
rect 503924 436624 503976 436640
rect 503716 436590 503740 436624
rect 503740 436590 503768 436624
rect 503820 436590 503840 436624
rect 503840 436590 503872 436624
rect 503924 436590 503940 436624
rect 503940 436590 503974 436624
rect 503974 436590 503976 436624
rect 503716 436588 503768 436590
rect 503820 436588 503872 436590
rect 503924 436588 503976 436590
rect 504028 436624 504080 436640
rect 504028 436590 504040 436624
rect 504040 436590 504074 436624
rect 504074 436590 504080 436624
rect 504028 436588 504080 436590
rect 504132 436624 504184 436640
rect 504132 436590 504140 436624
rect 504140 436590 504174 436624
rect 504174 436590 504184 436624
rect 504132 436588 504184 436590
rect 504236 436624 504288 436640
rect 504236 436590 504240 436624
rect 504240 436590 504274 436624
rect 504274 436590 504288 436624
rect 504236 436588 504288 436590
rect 503716 436524 503768 436536
rect 503820 436524 503872 436536
rect 503924 436524 503976 436536
rect 503716 436490 503740 436524
rect 503740 436490 503768 436524
rect 503820 436490 503840 436524
rect 503840 436490 503872 436524
rect 503924 436490 503940 436524
rect 503940 436490 503974 436524
rect 503974 436490 503976 436524
rect 503716 436484 503768 436490
rect 503820 436484 503872 436490
rect 503924 436484 503976 436490
rect 504028 436524 504080 436536
rect 504028 436490 504040 436524
rect 504040 436490 504074 436524
rect 504074 436490 504080 436524
rect 504028 436484 504080 436490
rect 504132 436524 504184 436536
rect 504132 436490 504140 436524
rect 504140 436490 504174 436524
rect 504174 436490 504184 436524
rect 504132 436484 504184 436490
rect 504236 436524 504288 436536
rect 504236 436490 504240 436524
rect 504240 436490 504274 436524
rect 504274 436490 504288 436524
rect 504236 436484 504288 436490
rect 503716 436424 503768 436432
rect 503820 436424 503872 436432
rect 503924 436424 503976 436432
rect 503716 436390 503740 436424
rect 503740 436390 503768 436424
rect 503820 436390 503840 436424
rect 503840 436390 503872 436424
rect 503924 436390 503940 436424
rect 503940 436390 503974 436424
rect 503974 436390 503976 436424
rect 503716 436380 503768 436390
rect 503820 436380 503872 436390
rect 503924 436380 503976 436390
rect 504028 436424 504080 436432
rect 504028 436390 504040 436424
rect 504040 436390 504074 436424
rect 504074 436390 504080 436424
rect 504028 436380 504080 436390
rect 504132 436424 504184 436432
rect 504132 436390 504140 436424
rect 504140 436390 504174 436424
rect 504174 436390 504184 436424
rect 504132 436380 504184 436390
rect 504236 436424 504288 436432
rect 504236 436390 504240 436424
rect 504240 436390 504274 436424
rect 504274 436390 504288 436424
rect 504236 436380 504288 436390
rect 503716 436324 503768 436328
rect 503820 436324 503872 436328
rect 503924 436324 503976 436328
rect 503716 436290 503740 436324
rect 503740 436290 503768 436324
rect 503820 436290 503840 436324
rect 503840 436290 503872 436324
rect 503924 436290 503940 436324
rect 503940 436290 503974 436324
rect 503974 436290 503976 436324
rect 503716 436276 503768 436290
rect 503820 436276 503872 436290
rect 503924 436276 503976 436290
rect 504028 436324 504080 436328
rect 504028 436290 504040 436324
rect 504040 436290 504074 436324
rect 504074 436290 504080 436324
rect 504028 436276 504080 436290
rect 504132 436324 504184 436328
rect 504132 436290 504140 436324
rect 504140 436290 504174 436324
rect 504174 436290 504184 436324
rect 504132 436276 504184 436290
rect 504236 436324 504288 436328
rect 504236 436290 504240 436324
rect 504240 436290 504274 436324
rect 504274 436290 504288 436324
rect 504236 436276 504288 436290
rect 508868 435536 508920 435560
rect 508972 435536 509024 435560
rect 509076 435536 509128 435560
rect 508868 435508 508892 435536
rect 508892 435508 508920 435536
rect 508972 435508 508992 435536
rect 508992 435508 509024 435536
rect 509076 435508 509092 435536
rect 509092 435508 509126 435536
rect 509126 435508 509128 435536
rect 509180 435536 509232 435560
rect 509180 435508 509192 435536
rect 509192 435508 509226 435536
rect 509226 435508 509232 435536
rect 509284 435536 509336 435560
rect 509284 435508 509292 435536
rect 509292 435508 509326 435536
rect 509326 435508 509336 435536
rect 509388 435536 509440 435560
rect 509388 435508 509392 435536
rect 509392 435508 509426 435536
rect 509426 435508 509440 435536
rect 508868 435436 508920 435456
rect 508972 435436 509024 435456
rect 509076 435436 509128 435456
rect 508868 435404 508892 435436
rect 508892 435404 508920 435436
rect 508972 435404 508992 435436
rect 508992 435404 509024 435436
rect 509076 435404 509092 435436
rect 509092 435404 509126 435436
rect 509126 435404 509128 435436
rect 509180 435436 509232 435456
rect 509180 435404 509192 435436
rect 509192 435404 509226 435436
rect 509226 435404 509232 435436
rect 509284 435436 509336 435456
rect 509284 435404 509292 435436
rect 509292 435404 509326 435436
rect 509326 435404 509336 435436
rect 509388 435436 509440 435456
rect 509388 435404 509392 435436
rect 509392 435404 509426 435436
rect 509426 435404 509440 435436
rect 508868 435336 508920 435352
rect 508972 435336 509024 435352
rect 509076 435336 509128 435352
rect 508868 435302 508892 435336
rect 508892 435302 508920 435336
rect 508972 435302 508992 435336
rect 508992 435302 509024 435336
rect 509076 435302 509092 435336
rect 509092 435302 509126 435336
rect 509126 435302 509128 435336
rect 508868 435300 508920 435302
rect 508972 435300 509024 435302
rect 509076 435300 509128 435302
rect 509180 435336 509232 435352
rect 509180 435302 509192 435336
rect 509192 435302 509226 435336
rect 509226 435302 509232 435336
rect 509180 435300 509232 435302
rect 509284 435336 509336 435352
rect 509284 435302 509292 435336
rect 509292 435302 509326 435336
rect 509326 435302 509336 435336
rect 509284 435300 509336 435302
rect 509388 435336 509440 435352
rect 509388 435302 509392 435336
rect 509392 435302 509426 435336
rect 509426 435302 509440 435336
rect 509388 435300 509440 435302
rect 508868 435236 508920 435248
rect 508972 435236 509024 435248
rect 509076 435236 509128 435248
rect 508868 435202 508892 435236
rect 508892 435202 508920 435236
rect 508972 435202 508992 435236
rect 508992 435202 509024 435236
rect 509076 435202 509092 435236
rect 509092 435202 509126 435236
rect 509126 435202 509128 435236
rect 508868 435196 508920 435202
rect 508972 435196 509024 435202
rect 509076 435196 509128 435202
rect 509180 435236 509232 435248
rect 509180 435202 509192 435236
rect 509192 435202 509226 435236
rect 509226 435202 509232 435236
rect 509180 435196 509232 435202
rect 509284 435236 509336 435248
rect 509284 435202 509292 435236
rect 509292 435202 509326 435236
rect 509326 435202 509336 435236
rect 509284 435196 509336 435202
rect 509388 435236 509440 435248
rect 509388 435202 509392 435236
rect 509392 435202 509426 435236
rect 509426 435202 509440 435236
rect 509388 435196 509440 435202
rect 508868 435136 508920 435144
rect 508972 435136 509024 435144
rect 509076 435136 509128 435144
rect 508868 435102 508892 435136
rect 508892 435102 508920 435136
rect 508972 435102 508992 435136
rect 508992 435102 509024 435136
rect 509076 435102 509092 435136
rect 509092 435102 509126 435136
rect 509126 435102 509128 435136
rect 508868 435092 508920 435102
rect 508972 435092 509024 435102
rect 509076 435092 509128 435102
rect 509180 435136 509232 435144
rect 509180 435102 509192 435136
rect 509192 435102 509226 435136
rect 509226 435102 509232 435136
rect 509180 435092 509232 435102
rect 509284 435136 509336 435144
rect 509284 435102 509292 435136
rect 509292 435102 509326 435136
rect 509326 435102 509336 435136
rect 509284 435092 509336 435102
rect 509388 435136 509440 435144
rect 509388 435102 509392 435136
rect 509392 435102 509426 435136
rect 509426 435102 509440 435136
rect 509388 435092 509440 435102
rect 508868 435036 508920 435040
rect 508972 435036 509024 435040
rect 509076 435036 509128 435040
rect 508868 435002 508892 435036
rect 508892 435002 508920 435036
rect 508972 435002 508992 435036
rect 508992 435002 509024 435036
rect 509076 435002 509092 435036
rect 509092 435002 509126 435036
rect 509126 435002 509128 435036
rect 508868 434988 508920 435002
rect 508972 434988 509024 435002
rect 509076 434988 509128 435002
rect 509180 435036 509232 435040
rect 509180 435002 509192 435036
rect 509192 435002 509226 435036
rect 509226 435002 509232 435036
rect 509180 434988 509232 435002
rect 509284 435036 509336 435040
rect 509284 435002 509292 435036
rect 509292 435002 509326 435036
rect 509326 435002 509336 435036
rect 509284 434988 509336 435002
rect 509388 435036 509440 435040
rect 509388 435002 509392 435036
rect 509392 435002 509426 435036
rect 509426 435002 509440 435036
rect 509388 434988 509440 435002
rect 527638 437440 527738 437540
rect 527862 437440 527962 437540
rect 528086 437440 528186 437540
rect 528310 437440 528410 437540
rect 528534 437440 528634 437540
rect 527638 437216 527738 437316
rect 527862 437216 527962 437316
rect 528086 437216 528186 437316
rect 528310 437216 528410 437316
rect 528534 437216 528634 437316
rect 527638 436992 527738 437092
rect 527862 436992 527962 437092
rect 528086 436992 528186 437092
rect 528310 436992 528410 437092
rect 528534 436992 528634 437092
rect 527638 436768 527738 436868
rect 527862 436768 527962 436868
rect 528086 436768 528186 436868
rect 528310 436768 528410 436868
rect 528534 436768 528634 436868
rect 527638 436544 527738 436644
rect 527862 436544 527962 436644
rect 528086 436544 528186 436644
rect 528310 436544 528410 436644
rect 528534 436544 528634 436644
rect 527638 436320 527738 436420
rect 527862 436320 527962 436420
rect 528086 436320 528186 436420
rect 528310 436320 528410 436420
rect 528534 436320 528634 436420
rect 527638 436096 527738 436196
rect 527862 436096 527962 436196
rect 528086 436096 528186 436196
rect 528310 436096 528410 436196
rect 528534 436096 528634 436196
rect 527638 435872 527738 435972
rect 527862 435872 527962 435972
rect 528086 435872 528186 435972
rect 528310 435872 528410 435972
rect 528534 435872 528634 435972
rect 527638 435648 527738 435748
rect 527862 435648 527962 435748
rect 528086 435648 528186 435748
rect 528310 435648 528410 435748
rect 528534 435648 528634 435748
rect 527638 435424 527738 435524
rect 527862 435424 527962 435524
rect 528086 435424 528186 435524
rect 528310 435424 528410 435524
rect 528534 435424 528634 435524
rect 527638 435200 527738 435300
rect 527862 435200 527962 435300
rect 528086 435200 528186 435300
rect 528310 435200 528410 435300
rect 528534 435200 528634 435300
rect 527638 434976 527738 435076
rect 527862 434976 527962 435076
rect 528086 434976 528186 435076
rect 528310 434976 528410 435076
rect 528534 434976 528634 435076
rect 527638 434752 527738 434852
rect 527862 434752 527962 434852
rect 528086 434752 528186 434852
rect 528310 434752 528410 434852
rect 528534 434752 528634 434852
rect 527638 434528 527738 434628
rect 527862 434528 527962 434628
rect 528086 434528 528186 434628
rect 528310 434528 528410 434628
rect 528534 434528 528634 434628
rect 527638 434304 527738 434404
rect 527862 434304 527962 434404
rect 528086 434304 528186 434404
rect 528310 434304 528410 434404
rect 528534 434304 528634 434404
rect 527638 434080 527738 434180
rect 527862 434080 527962 434180
rect 528086 434080 528186 434180
rect 528310 434080 528410 434180
rect 528534 434080 528634 434180
rect 527638 433856 527738 433956
rect 527862 433856 527962 433956
rect 528086 433856 528186 433956
rect 528310 433856 528410 433956
rect 528534 433856 528634 433956
rect 527638 433632 527738 433732
rect 527862 433632 527962 433732
rect 528086 433632 528186 433732
rect 528310 433632 528410 433732
rect 528534 433632 528634 433732
rect 527638 433408 527738 433508
rect 527862 433408 527962 433508
rect 528086 433408 528186 433508
rect 528310 433408 528410 433508
rect 528534 433408 528634 433508
rect 527638 433184 527738 433284
rect 527862 433184 527962 433284
rect 528086 433184 528186 433284
rect 528310 433184 528410 433284
rect 528534 433184 528634 433284
rect 527638 432960 527738 433060
rect 527862 432960 527962 433060
rect 528086 432960 528186 433060
rect 528310 432960 528410 433060
rect 528534 432960 528634 433060
rect 527638 432736 527738 432836
rect 527862 432736 527962 432836
rect 528086 432736 528186 432836
rect 528310 432736 528410 432836
rect 528534 432736 528634 432836
rect 527638 432512 527738 432612
rect 527862 432512 527962 432612
rect 528086 432512 528186 432612
rect 528310 432512 528410 432612
rect 528534 432512 528634 432612
rect 500418 432064 500518 432164
rect 500642 432064 500742 432164
rect 500866 432064 500966 432164
rect 501090 432064 501190 432164
rect 501314 432064 501414 432164
rect 500418 431840 500518 431940
rect 500642 431840 500742 431940
rect 500866 431840 500966 431940
rect 501090 431840 501190 431940
rect 501314 431840 501414 431940
rect 500418 431616 500518 431716
rect 500642 431616 500742 431716
rect 500866 431616 500966 431716
rect 501090 431616 501190 431716
rect 501314 431616 501414 431716
rect 500418 431392 500518 431492
rect 500642 431392 500742 431492
rect 500866 431392 500966 431492
rect 501090 431392 501190 431492
rect 501314 431392 501414 431492
rect 500418 431168 500518 431268
rect 500642 431168 500742 431268
rect 500866 431168 500966 431268
rect 501090 431168 501190 431268
rect 501314 431168 501414 431268
rect 527638 432288 527738 432388
rect 527862 432288 527962 432388
rect 528086 432288 528186 432388
rect 528310 432288 528410 432388
rect 528534 432288 528634 432388
rect 527638 432064 527738 432164
rect 527862 432064 527962 432164
rect 528086 432064 528186 432164
rect 528310 432064 528410 432164
rect 528534 432064 528634 432164
rect 527638 431840 527738 431940
rect 527862 431840 527962 431940
rect 528086 431840 528186 431940
rect 528310 431840 528410 431940
rect 528534 431840 528634 431940
rect 527638 431616 527738 431716
rect 527862 431616 527962 431716
rect 528086 431616 528186 431716
rect 528310 431616 528410 431716
rect 528534 431616 528634 431716
rect 527638 431392 527738 431492
rect 527862 431392 527962 431492
rect 528086 431392 528186 431492
rect 528310 431392 528410 431492
rect 528534 431392 528634 431492
rect 527638 431168 527738 431268
rect 527862 431168 527962 431268
rect 528086 431168 528186 431268
rect 528310 431168 528410 431268
rect 528534 431168 528634 431268
rect 500418 430944 500518 431044
rect 500642 430944 500742 431044
rect 500866 430944 500966 431044
rect 501090 430944 501190 431044
rect 501314 430944 501414 431044
rect 503920 430926 504020 431026
rect 504144 430926 504244 431026
rect 504368 430926 504468 431026
rect 504592 430926 504692 431026
rect 504816 430926 504916 431026
rect 505040 430926 505140 431026
rect 505264 430926 505364 431026
rect 505488 430926 505588 431026
rect 505712 430926 505812 431026
rect 505936 430926 506036 431026
rect 506160 430926 506260 431026
rect 506384 430926 506484 431026
rect 506608 430926 506708 431026
rect 506832 430926 506932 431026
rect 507056 430926 507156 431026
rect 507280 430926 507380 431026
rect 507504 430926 507604 431026
rect 507728 430926 507828 431026
rect 507952 430926 508052 431026
rect 508176 430926 508276 431026
rect 508400 430926 508500 431026
rect 508624 430926 508724 431026
rect 508848 430926 508948 431026
rect 509072 430926 509172 431026
rect 509296 430926 509396 431026
rect 509520 430926 509620 431026
rect 509744 430926 509844 431026
rect 509968 430926 510068 431026
rect 510192 430926 510292 431026
rect 510416 430926 510516 431026
rect 503920 430702 504020 430802
rect 504144 430702 504244 430802
rect 504368 430702 504468 430802
rect 504592 430702 504692 430802
rect 504816 430702 504916 430802
rect 505040 430702 505140 430802
rect 505264 430702 505364 430802
rect 505488 430702 505588 430802
rect 505712 430702 505812 430802
rect 505936 430702 506036 430802
rect 506160 430702 506260 430802
rect 506384 430702 506484 430802
rect 506608 430702 506708 430802
rect 506832 430702 506932 430802
rect 507056 430702 507156 430802
rect 507280 430702 507380 430802
rect 507504 430702 507604 430802
rect 507728 430702 507828 430802
rect 507952 430702 508052 430802
rect 508176 430702 508276 430802
rect 508400 430702 508500 430802
rect 508624 430702 508724 430802
rect 508848 430702 508948 430802
rect 509072 430702 509172 430802
rect 509296 430702 509396 430802
rect 509520 430702 509620 430802
rect 509744 430702 509844 430802
rect 509968 430702 510068 430802
rect 510192 430702 510292 430802
rect 510416 430702 510516 430802
rect 503920 430478 504020 430578
rect 504144 430478 504244 430578
rect 504368 430478 504468 430578
rect 504592 430478 504692 430578
rect 504816 430478 504916 430578
rect 505040 430478 505140 430578
rect 505264 430478 505364 430578
rect 505488 430478 505588 430578
rect 505712 430478 505812 430578
rect 505936 430478 506036 430578
rect 506160 430478 506260 430578
rect 506384 430478 506484 430578
rect 506608 430478 506708 430578
rect 506832 430478 506932 430578
rect 507056 430478 507156 430578
rect 507280 430478 507380 430578
rect 507504 430478 507604 430578
rect 507728 430478 507828 430578
rect 507952 430478 508052 430578
rect 508176 430478 508276 430578
rect 508400 430478 508500 430578
rect 508624 430478 508724 430578
rect 508848 430478 508948 430578
rect 509072 430478 509172 430578
rect 509296 430478 509396 430578
rect 509520 430478 509620 430578
rect 509744 430478 509844 430578
rect 509968 430478 510068 430578
rect 510192 430478 510292 430578
rect 510416 430478 510516 430578
rect 503920 430254 504020 430354
rect 504144 430254 504244 430354
rect 504368 430254 504468 430354
rect 504592 430254 504692 430354
rect 504816 430254 504916 430354
rect 505040 430254 505140 430354
rect 505264 430254 505364 430354
rect 505488 430254 505588 430354
rect 505712 430254 505812 430354
rect 505936 430254 506036 430354
rect 506160 430254 506260 430354
rect 506384 430254 506484 430354
rect 506608 430254 506708 430354
rect 506832 430254 506932 430354
rect 507056 430254 507156 430354
rect 507280 430254 507380 430354
rect 507504 430254 507604 430354
rect 507728 430254 507828 430354
rect 507952 430254 508052 430354
rect 508176 430254 508276 430354
rect 508400 430254 508500 430354
rect 508624 430254 508724 430354
rect 508848 430254 508948 430354
rect 509072 430254 509172 430354
rect 509296 430254 509396 430354
rect 509520 430254 509620 430354
rect 509744 430254 509844 430354
rect 509968 430254 510068 430354
rect 510192 430254 510292 430354
rect 510416 430254 510516 430354
rect 503920 430030 504020 430130
rect 504144 430030 504244 430130
rect 504368 430030 504468 430130
rect 504592 430030 504692 430130
rect 504816 430030 504916 430130
rect 505040 430030 505140 430130
rect 505264 430030 505364 430130
rect 505488 430030 505588 430130
rect 505712 430030 505812 430130
rect 505936 430030 506036 430130
rect 506160 430030 506260 430130
rect 506384 430030 506484 430130
rect 506608 430030 506708 430130
rect 506832 430030 506932 430130
rect 507056 430030 507156 430130
rect 507280 430030 507380 430130
rect 507504 430030 507604 430130
rect 507728 430030 507828 430130
rect 507952 430030 508052 430130
rect 508176 430030 508276 430130
rect 508400 430030 508500 430130
rect 508624 430030 508724 430130
rect 508848 430030 508948 430130
rect 509072 430030 509172 430130
rect 509296 430030 509396 430130
rect 509520 430030 509620 430130
rect 509744 430030 509844 430130
rect 509968 430030 510068 430130
rect 510192 430030 510292 430130
rect 510416 430030 510516 430130
rect 517320 430926 517420 431026
rect 517544 430926 517644 431026
rect 517768 430926 517868 431026
rect 517992 430926 518092 431026
rect 518216 430926 518316 431026
rect 518440 430926 518540 431026
rect 518664 430926 518764 431026
rect 518888 430926 518988 431026
rect 519112 430926 519212 431026
rect 519336 430926 519436 431026
rect 519560 430926 519660 431026
rect 519784 430926 519884 431026
rect 520008 430926 520108 431026
rect 520232 430926 520332 431026
rect 520456 430926 520556 431026
rect 520680 430926 520780 431026
rect 520904 430926 521004 431026
rect 521128 430926 521228 431026
rect 521352 430926 521452 431026
rect 521576 430926 521676 431026
rect 521800 430926 521900 431026
rect 522024 430926 522124 431026
rect 522248 430926 522348 431026
rect 522472 430926 522572 431026
rect 522696 430926 522796 431026
rect 522920 430926 523020 431026
rect 523144 430926 523244 431026
rect 523368 430926 523468 431026
rect 523592 430926 523692 431026
rect 523816 430926 523916 431026
rect 527638 430944 527738 431044
rect 527862 430944 527962 431044
rect 528086 430944 528186 431044
rect 528310 430944 528410 431044
rect 528534 430944 528634 431044
rect 517320 430702 517420 430802
rect 517544 430702 517644 430802
rect 517768 430702 517868 430802
rect 517992 430702 518092 430802
rect 518216 430702 518316 430802
rect 518440 430702 518540 430802
rect 518664 430702 518764 430802
rect 518888 430702 518988 430802
rect 519112 430702 519212 430802
rect 519336 430702 519436 430802
rect 519560 430702 519660 430802
rect 519784 430702 519884 430802
rect 520008 430702 520108 430802
rect 520232 430702 520332 430802
rect 520456 430702 520556 430802
rect 520680 430702 520780 430802
rect 520904 430702 521004 430802
rect 521128 430702 521228 430802
rect 521352 430702 521452 430802
rect 521576 430702 521676 430802
rect 521800 430702 521900 430802
rect 522024 430702 522124 430802
rect 522248 430702 522348 430802
rect 522472 430702 522572 430802
rect 522696 430702 522796 430802
rect 522920 430702 523020 430802
rect 523144 430702 523244 430802
rect 523368 430702 523468 430802
rect 523592 430702 523692 430802
rect 523816 430702 523916 430802
rect 517320 430478 517420 430578
rect 517544 430478 517644 430578
rect 517768 430478 517868 430578
rect 517992 430478 518092 430578
rect 518216 430478 518316 430578
rect 518440 430478 518540 430578
rect 518664 430478 518764 430578
rect 518888 430478 518988 430578
rect 519112 430478 519212 430578
rect 519336 430478 519436 430578
rect 519560 430478 519660 430578
rect 519784 430478 519884 430578
rect 520008 430478 520108 430578
rect 520232 430478 520332 430578
rect 520456 430478 520556 430578
rect 520680 430478 520780 430578
rect 520904 430478 521004 430578
rect 521128 430478 521228 430578
rect 521352 430478 521452 430578
rect 521576 430478 521676 430578
rect 521800 430478 521900 430578
rect 522024 430478 522124 430578
rect 522248 430478 522348 430578
rect 522472 430478 522572 430578
rect 522696 430478 522796 430578
rect 522920 430478 523020 430578
rect 523144 430478 523244 430578
rect 523368 430478 523468 430578
rect 523592 430478 523692 430578
rect 523816 430478 523916 430578
rect 517320 430254 517420 430354
rect 517544 430254 517644 430354
rect 517768 430254 517868 430354
rect 517992 430254 518092 430354
rect 518216 430254 518316 430354
rect 518440 430254 518540 430354
rect 518664 430254 518764 430354
rect 518888 430254 518988 430354
rect 519112 430254 519212 430354
rect 519336 430254 519436 430354
rect 519560 430254 519660 430354
rect 519784 430254 519884 430354
rect 520008 430254 520108 430354
rect 520232 430254 520332 430354
rect 520456 430254 520556 430354
rect 520680 430254 520780 430354
rect 520904 430254 521004 430354
rect 521128 430254 521228 430354
rect 521352 430254 521452 430354
rect 521576 430254 521676 430354
rect 521800 430254 521900 430354
rect 522024 430254 522124 430354
rect 522248 430254 522348 430354
rect 522472 430254 522572 430354
rect 522696 430254 522796 430354
rect 522920 430254 523020 430354
rect 523144 430254 523244 430354
rect 523368 430254 523468 430354
rect 523592 430254 523692 430354
rect 523816 430254 523916 430354
rect 517320 430030 517420 430130
rect 517544 430030 517644 430130
rect 517768 430030 517868 430130
rect 517992 430030 518092 430130
rect 518216 430030 518316 430130
rect 518440 430030 518540 430130
rect 518664 430030 518764 430130
rect 518888 430030 518988 430130
rect 519112 430030 519212 430130
rect 519336 430030 519436 430130
rect 519560 430030 519660 430130
rect 519784 430030 519884 430130
rect 520008 430030 520108 430130
rect 520232 430030 520332 430130
rect 520456 430030 520556 430130
rect 520680 430030 520780 430130
rect 520904 430030 521004 430130
rect 521128 430030 521228 430130
rect 521352 430030 521452 430130
rect 521576 430030 521676 430130
rect 521800 430030 521900 430130
rect 522024 430030 522124 430130
rect 522248 430030 522348 430130
rect 522472 430030 522572 430130
rect 522696 430030 522796 430130
rect 522920 430030 523020 430130
rect 523144 430030 523244 430130
rect 523368 430030 523468 430130
rect 523592 430030 523692 430130
rect 523816 430030 523916 430130
<< metal2 >>
rect 562380 495742 567480 495822
rect 562380 495662 562480 495742
rect 562560 495662 562640 495742
rect 562720 495662 562800 495742
rect 562880 495662 562960 495742
rect 563040 495662 563120 495742
rect 563200 495662 563280 495742
rect 563360 495662 563440 495742
rect 563520 495662 563600 495742
rect 563680 495662 563760 495742
rect 563840 495662 563920 495742
rect 564000 495662 564080 495742
rect 564160 495662 564240 495742
rect 564320 495662 564400 495742
rect 564480 495662 564560 495742
rect 564640 495662 564720 495742
rect 564800 495662 564880 495742
rect 564960 495662 565040 495742
rect 565120 495662 565200 495742
rect 565280 495662 565360 495742
rect 565440 495662 565520 495742
rect 565600 495662 565680 495742
rect 565760 495662 565840 495742
rect 565920 495662 566000 495742
rect 566080 495662 566160 495742
rect 566240 495662 566320 495742
rect 566400 495662 566480 495742
rect 566560 495662 566640 495742
rect 566720 495662 566800 495742
rect 566880 495662 566960 495742
rect 567040 495662 567120 495742
rect 567200 495662 567280 495742
rect 567360 495662 567480 495742
rect 562380 495582 567480 495662
rect 562380 495502 562480 495582
rect 562560 495502 562640 495582
rect 562720 495502 562800 495582
rect 562880 495502 562960 495582
rect 563040 495502 563120 495582
rect 563200 495502 563280 495582
rect 563360 495502 563440 495582
rect 563520 495502 563600 495582
rect 563680 495502 563760 495582
rect 563840 495502 563920 495582
rect 564000 495502 564080 495582
rect 564160 495502 564240 495582
rect 564320 495502 564400 495582
rect 564480 495502 564560 495582
rect 564640 495502 564720 495582
rect 564800 495502 564880 495582
rect 564960 495502 565040 495582
rect 565120 495502 565200 495582
rect 565280 495502 565360 495582
rect 565440 495502 565520 495582
rect 565600 495502 565680 495582
rect 565760 495502 565840 495582
rect 565920 495502 566000 495582
rect 566080 495502 566160 495582
rect 566240 495502 566320 495582
rect 566400 495502 566480 495582
rect 566560 495502 566640 495582
rect 566720 495502 566800 495582
rect 566880 495502 566960 495582
rect 567040 495502 567120 495582
rect 567200 495502 567280 495582
rect 567360 495502 567480 495582
rect 562380 495462 567480 495502
rect 572540 495742 577640 495822
rect 572540 495662 572640 495742
rect 572720 495662 572800 495742
rect 572880 495662 572960 495742
rect 573040 495662 573120 495742
rect 573200 495662 573280 495742
rect 573360 495662 573440 495742
rect 573520 495662 573600 495742
rect 573680 495662 573760 495742
rect 573840 495662 573920 495742
rect 574000 495662 574080 495742
rect 574160 495662 574240 495742
rect 574320 495662 574400 495742
rect 574480 495662 574560 495742
rect 574640 495662 574720 495742
rect 574800 495662 574880 495742
rect 574960 495662 575040 495742
rect 575120 495662 575200 495742
rect 575280 495662 575360 495742
rect 575440 495662 575520 495742
rect 575600 495662 575680 495742
rect 575760 495662 575840 495742
rect 575920 495662 576000 495742
rect 576080 495662 576160 495742
rect 576240 495662 576320 495742
rect 576400 495662 576480 495742
rect 576560 495662 576640 495742
rect 576720 495662 576800 495742
rect 576880 495662 576960 495742
rect 577040 495662 577120 495742
rect 577200 495662 577280 495742
rect 577360 495662 577440 495742
rect 577520 495662 577640 495742
rect 572540 495582 577640 495662
rect 572540 495502 572640 495582
rect 572720 495502 572800 495582
rect 572880 495502 572960 495582
rect 573040 495502 573120 495582
rect 573200 495502 573280 495582
rect 573360 495502 573440 495582
rect 573520 495502 573600 495582
rect 573680 495502 573760 495582
rect 573840 495502 573920 495582
rect 574000 495502 574080 495582
rect 574160 495502 574240 495582
rect 574320 495502 574400 495582
rect 574480 495502 574560 495582
rect 574640 495502 574720 495582
rect 574800 495502 574880 495582
rect 574960 495502 575040 495582
rect 575120 495502 575200 495582
rect 575280 495502 575360 495582
rect 575440 495502 575520 495582
rect 575600 495502 575680 495582
rect 575760 495502 575840 495582
rect 575920 495502 576000 495582
rect 576080 495502 576160 495582
rect 576240 495502 576320 495582
rect 576400 495502 576480 495582
rect 576560 495502 576640 495582
rect 576720 495502 576800 495582
rect 576880 495502 576960 495582
rect 577040 495502 577120 495582
rect 577200 495502 577280 495582
rect 577360 495502 577440 495582
rect 577520 495502 577640 495582
rect 572540 495462 577640 495502
rect 562102 494221 567622 494281
rect 562102 494161 562222 494221
rect 562282 494161 562342 494221
rect 562402 494161 562462 494221
rect 562522 494161 562582 494221
rect 562642 494161 562702 494221
rect 562762 494161 562822 494221
rect 562882 494161 562942 494221
rect 563002 494161 563062 494221
rect 563122 494161 563182 494221
rect 563242 494161 563302 494221
rect 563362 494161 563422 494221
rect 563482 494161 563542 494221
rect 563602 494161 563662 494221
rect 563722 494161 563782 494221
rect 563842 494161 563902 494221
rect 563962 494161 564022 494221
rect 564082 494161 564142 494221
rect 564202 494161 564262 494221
rect 564322 494161 564382 494221
rect 564442 494161 564502 494221
rect 564562 494161 564622 494221
rect 564682 494161 564742 494221
rect 564802 494161 564862 494221
rect 564922 494161 564982 494221
rect 565042 494161 565102 494221
rect 565162 494161 565222 494221
rect 565282 494161 565342 494221
rect 565402 494161 565462 494221
rect 565522 494161 565582 494221
rect 565642 494161 565702 494221
rect 565762 494161 565822 494221
rect 565882 494161 565942 494221
rect 566002 494161 566062 494221
rect 566122 494161 566182 494221
rect 566242 494161 566302 494221
rect 566362 494161 566422 494221
rect 566482 494161 566542 494221
rect 566602 494161 566662 494221
rect 566722 494161 566782 494221
rect 566842 494161 566902 494221
rect 566962 494161 567022 494221
rect 567082 494161 567142 494221
rect 567202 494161 567262 494221
rect 567322 494161 567382 494221
rect 567442 494161 567502 494221
rect 567562 494161 567622 494221
rect 562102 494101 567622 494161
rect 562102 494041 562222 494101
rect 562282 494041 562342 494101
rect 562402 494041 562462 494101
rect 562522 494041 562582 494101
rect 562642 494041 562702 494101
rect 562762 494041 562822 494101
rect 562882 494041 562942 494101
rect 563002 494041 563062 494101
rect 563122 494041 563182 494101
rect 563242 494041 563302 494101
rect 563362 494041 563422 494101
rect 563482 494041 563542 494101
rect 563602 494041 563662 494101
rect 563722 494041 563782 494101
rect 563842 494041 563902 494101
rect 563962 494041 564022 494101
rect 564082 494041 564142 494101
rect 564202 494041 564262 494101
rect 564322 494041 564382 494101
rect 564442 494041 564502 494101
rect 564562 494041 564622 494101
rect 564682 494041 564742 494101
rect 564802 494041 564862 494101
rect 564922 494041 564982 494101
rect 565042 494041 565102 494101
rect 565162 494041 565222 494101
rect 565282 494041 565342 494101
rect 565402 494041 565462 494101
rect 565522 494041 565582 494101
rect 565642 494041 565702 494101
rect 565762 494041 565822 494101
rect 565882 494041 565942 494101
rect 566002 494041 566062 494101
rect 566122 494041 566182 494101
rect 566242 494041 566302 494101
rect 566362 494041 566422 494101
rect 566482 494041 566542 494101
rect 566602 494041 566662 494101
rect 566722 494041 566782 494101
rect 566842 494041 566902 494101
rect 566962 494041 567022 494101
rect 567082 494041 567142 494101
rect 567202 494041 567262 494101
rect 567322 494041 567382 494101
rect 567442 494041 567502 494101
rect 567562 494041 567622 494101
rect 562102 493981 567622 494041
rect 572272 494236 577792 494296
rect 572272 494176 572332 494236
rect 572392 494176 572452 494236
rect 572512 494176 572572 494236
rect 572632 494176 572692 494236
rect 572752 494176 572812 494236
rect 572872 494176 572932 494236
rect 572992 494176 573052 494236
rect 573112 494176 573172 494236
rect 573232 494176 573292 494236
rect 573352 494176 573412 494236
rect 573472 494176 573532 494236
rect 573592 494176 573652 494236
rect 573712 494176 573772 494236
rect 573832 494176 573892 494236
rect 573952 494176 574012 494236
rect 574072 494176 574132 494236
rect 574192 494176 574252 494236
rect 574312 494176 574372 494236
rect 574432 494176 574492 494236
rect 574552 494176 574612 494236
rect 574672 494176 574732 494236
rect 574792 494176 574852 494236
rect 574912 494176 574972 494236
rect 575032 494176 575092 494236
rect 575152 494176 575212 494236
rect 575272 494176 575332 494236
rect 575392 494176 575452 494236
rect 575512 494176 575572 494236
rect 575632 494176 575692 494236
rect 575752 494176 575812 494236
rect 575872 494176 575932 494236
rect 575992 494176 576052 494236
rect 576112 494176 576172 494236
rect 576232 494176 576292 494236
rect 576352 494176 576412 494236
rect 576472 494176 576532 494236
rect 576592 494176 576652 494236
rect 576712 494176 576772 494236
rect 576832 494176 576892 494236
rect 576952 494176 577012 494236
rect 577072 494176 577132 494236
rect 577192 494176 577252 494236
rect 577312 494176 577372 494236
rect 577432 494176 577492 494236
rect 577552 494176 577612 494236
rect 577672 494176 577792 494236
rect 572272 494116 577792 494176
rect 572272 494056 572332 494116
rect 572392 494056 572452 494116
rect 572512 494056 572572 494116
rect 572632 494056 572692 494116
rect 572752 494056 572812 494116
rect 572872 494056 572932 494116
rect 572992 494056 573052 494116
rect 573112 494056 573172 494116
rect 573232 494056 573292 494116
rect 573352 494056 573412 494116
rect 573472 494056 573532 494116
rect 573592 494056 573652 494116
rect 573712 494056 573772 494116
rect 573832 494056 573892 494116
rect 573952 494056 574012 494116
rect 574072 494056 574132 494116
rect 574192 494056 574252 494116
rect 574312 494056 574372 494116
rect 574432 494056 574492 494116
rect 574552 494056 574612 494116
rect 574672 494056 574732 494116
rect 574792 494056 574852 494116
rect 574912 494056 574972 494116
rect 575032 494056 575092 494116
rect 575152 494056 575212 494116
rect 575272 494056 575332 494116
rect 575392 494056 575452 494116
rect 575512 494056 575572 494116
rect 575632 494056 575692 494116
rect 575752 494056 575812 494116
rect 575872 494056 575932 494116
rect 575992 494056 576052 494116
rect 576112 494056 576172 494116
rect 576232 494056 576292 494116
rect 576352 494056 576412 494116
rect 576472 494056 576532 494116
rect 576592 494056 576652 494116
rect 576712 494056 576772 494116
rect 576832 494056 576892 494116
rect 576952 494056 577012 494116
rect 577072 494056 577132 494116
rect 577192 494056 577252 494116
rect 577312 494056 577372 494116
rect 577432 494056 577492 494116
rect 577552 494056 577612 494116
rect 577672 494056 577792 494116
rect 572272 493996 577792 494056
rect 503900 475306 510526 475336
rect 503900 475206 503920 475306
rect 504020 475206 504144 475306
rect 504244 475206 504368 475306
rect 504468 475206 504592 475306
rect 504692 475206 504816 475306
rect 504916 475206 505040 475306
rect 505140 475206 505264 475306
rect 505364 475206 505488 475306
rect 505588 475206 505712 475306
rect 505812 475206 505936 475306
rect 506036 475206 506160 475306
rect 506260 475206 506384 475306
rect 506484 475206 506608 475306
rect 506708 475206 506832 475306
rect 506932 475206 507056 475306
rect 507156 475206 507280 475306
rect 507380 475206 507504 475306
rect 507604 475206 507728 475306
rect 507828 475206 507952 475306
rect 508052 475206 508176 475306
rect 508276 475206 508400 475306
rect 508500 475206 508624 475306
rect 508724 475206 508848 475306
rect 508948 475206 509072 475306
rect 509172 475206 509296 475306
rect 509396 475206 509520 475306
rect 509620 475206 509744 475306
rect 509844 475206 509968 475306
rect 510068 475206 510192 475306
rect 510292 475206 510416 475306
rect 510516 475206 510526 475306
rect 503900 475082 510526 475206
rect 503900 474982 503920 475082
rect 504020 474982 504144 475082
rect 504244 474982 504368 475082
rect 504468 474982 504592 475082
rect 504692 474982 504816 475082
rect 504916 474982 505040 475082
rect 505140 474982 505264 475082
rect 505364 474982 505488 475082
rect 505588 474982 505712 475082
rect 505812 474982 505936 475082
rect 506036 474982 506160 475082
rect 506260 474982 506384 475082
rect 506484 474982 506608 475082
rect 506708 474982 506832 475082
rect 506932 474982 507056 475082
rect 507156 474982 507280 475082
rect 507380 474982 507504 475082
rect 507604 474982 507728 475082
rect 507828 474982 507952 475082
rect 508052 474982 508176 475082
rect 508276 474982 508400 475082
rect 508500 474982 508624 475082
rect 508724 474982 508848 475082
rect 508948 474982 509072 475082
rect 509172 474982 509296 475082
rect 509396 474982 509520 475082
rect 509620 474982 509744 475082
rect 509844 474982 509968 475082
rect 510068 474982 510192 475082
rect 510292 474982 510416 475082
rect 510516 474982 510526 475082
rect 503900 474858 510526 474982
rect 503900 474758 503920 474858
rect 504020 474758 504144 474858
rect 504244 474758 504368 474858
rect 504468 474758 504592 474858
rect 504692 474758 504816 474858
rect 504916 474758 505040 474858
rect 505140 474758 505264 474858
rect 505364 474758 505488 474858
rect 505588 474758 505712 474858
rect 505812 474758 505936 474858
rect 506036 474758 506160 474858
rect 506260 474758 506384 474858
rect 506484 474758 506608 474858
rect 506708 474758 506832 474858
rect 506932 474758 507056 474858
rect 507156 474758 507280 474858
rect 507380 474758 507504 474858
rect 507604 474758 507728 474858
rect 507828 474758 507952 474858
rect 508052 474758 508176 474858
rect 508276 474758 508400 474858
rect 508500 474758 508624 474858
rect 508724 474758 508848 474858
rect 508948 474758 509072 474858
rect 509172 474758 509296 474858
rect 509396 474758 509520 474858
rect 509620 474758 509744 474858
rect 509844 474758 509968 474858
rect 510068 474758 510192 474858
rect 510292 474758 510416 474858
rect 510516 474758 510526 474858
rect 503900 474634 510526 474758
rect 503900 474534 503920 474634
rect 504020 474534 504144 474634
rect 504244 474534 504368 474634
rect 504468 474534 504592 474634
rect 504692 474534 504816 474634
rect 504916 474534 505040 474634
rect 505140 474534 505264 474634
rect 505364 474534 505488 474634
rect 505588 474534 505712 474634
rect 505812 474534 505936 474634
rect 506036 474534 506160 474634
rect 506260 474534 506384 474634
rect 506484 474534 506608 474634
rect 506708 474534 506832 474634
rect 506932 474534 507056 474634
rect 507156 474534 507280 474634
rect 507380 474534 507504 474634
rect 507604 474534 507728 474634
rect 507828 474534 507952 474634
rect 508052 474534 508176 474634
rect 508276 474534 508400 474634
rect 508500 474534 508624 474634
rect 508724 474534 508848 474634
rect 508948 474534 509072 474634
rect 509172 474534 509296 474634
rect 509396 474534 509520 474634
rect 509620 474534 509744 474634
rect 509844 474534 509968 474634
rect 510068 474534 510192 474634
rect 510292 474534 510416 474634
rect 510516 474534 510526 474634
rect 503900 474410 510526 474534
rect 500364 474280 501424 474320
rect 500364 474180 500398 474280
rect 500498 474180 500622 474280
rect 500722 474180 500846 474280
rect 500946 474180 501070 474280
rect 501170 474180 501294 474280
rect 501394 474180 501424 474280
rect 503900 474310 503920 474410
rect 504020 474310 504144 474410
rect 504244 474310 504368 474410
rect 504468 474310 504592 474410
rect 504692 474310 504816 474410
rect 504916 474310 505040 474410
rect 505140 474310 505264 474410
rect 505364 474310 505488 474410
rect 505588 474310 505712 474410
rect 505812 474310 505936 474410
rect 506036 474310 506160 474410
rect 506260 474310 506384 474410
rect 506484 474310 506608 474410
rect 506708 474310 506832 474410
rect 506932 474310 507056 474410
rect 507156 474310 507280 474410
rect 507380 474310 507504 474410
rect 507604 474310 507728 474410
rect 507828 474310 507952 474410
rect 508052 474310 508176 474410
rect 508276 474310 508400 474410
rect 508500 474310 508624 474410
rect 508724 474310 508848 474410
rect 508948 474310 509072 474410
rect 509172 474310 509296 474410
rect 509396 474310 509520 474410
rect 509620 474310 509744 474410
rect 509844 474310 509968 474410
rect 510068 474310 510192 474410
rect 510292 474310 510416 474410
rect 510516 474310 510526 474410
rect 503900 474278 510526 474310
rect 517280 475306 523940 475336
rect 517280 475206 517320 475306
rect 517420 475206 517544 475306
rect 517644 475206 517768 475306
rect 517868 475206 517992 475306
rect 518092 475206 518216 475306
rect 518316 475206 518440 475306
rect 518540 475206 518664 475306
rect 518764 475206 518888 475306
rect 518988 475206 519112 475306
rect 519212 475206 519336 475306
rect 519436 475206 519560 475306
rect 519660 475206 519784 475306
rect 519884 475206 520008 475306
rect 520108 475206 520232 475306
rect 520332 475206 520456 475306
rect 520556 475206 520680 475306
rect 520780 475206 520904 475306
rect 521004 475206 521128 475306
rect 521228 475206 521352 475306
rect 521452 475206 521576 475306
rect 521676 475206 521800 475306
rect 521900 475206 522024 475306
rect 522124 475206 522248 475306
rect 522348 475206 522472 475306
rect 522572 475206 522696 475306
rect 522796 475206 522920 475306
rect 523020 475206 523144 475306
rect 523244 475206 523368 475306
rect 523468 475206 523592 475306
rect 523692 475206 523816 475306
rect 523916 475206 523940 475306
rect 517280 475082 523940 475206
rect 517280 474982 517320 475082
rect 517420 474982 517544 475082
rect 517644 474982 517768 475082
rect 517868 474982 517992 475082
rect 518092 474982 518216 475082
rect 518316 474982 518440 475082
rect 518540 474982 518664 475082
rect 518764 474982 518888 475082
rect 518988 474982 519112 475082
rect 519212 474982 519336 475082
rect 519436 474982 519560 475082
rect 519660 474982 519784 475082
rect 519884 474982 520008 475082
rect 520108 474982 520232 475082
rect 520332 474982 520456 475082
rect 520556 474982 520680 475082
rect 520780 474982 520904 475082
rect 521004 474982 521128 475082
rect 521228 474982 521352 475082
rect 521452 474982 521576 475082
rect 521676 474982 521800 475082
rect 521900 474982 522024 475082
rect 522124 474982 522248 475082
rect 522348 474982 522472 475082
rect 522572 474982 522696 475082
rect 522796 474982 522920 475082
rect 523020 474982 523144 475082
rect 523244 474982 523368 475082
rect 523468 474982 523592 475082
rect 523692 474982 523816 475082
rect 523916 474982 523940 475082
rect 517280 474858 523940 474982
rect 517280 474758 517320 474858
rect 517420 474758 517544 474858
rect 517644 474758 517768 474858
rect 517868 474758 517992 474858
rect 518092 474758 518216 474858
rect 518316 474758 518440 474858
rect 518540 474758 518664 474858
rect 518764 474758 518888 474858
rect 518988 474758 519112 474858
rect 519212 474758 519336 474858
rect 519436 474758 519560 474858
rect 519660 474758 519784 474858
rect 519884 474758 520008 474858
rect 520108 474758 520232 474858
rect 520332 474758 520456 474858
rect 520556 474758 520680 474858
rect 520780 474758 520904 474858
rect 521004 474758 521128 474858
rect 521228 474758 521352 474858
rect 521452 474758 521576 474858
rect 521676 474758 521800 474858
rect 521900 474758 522024 474858
rect 522124 474758 522248 474858
rect 522348 474758 522472 474858
rect 522572 474758 522696 474858
rect 522796 474758 522920 474858
rect 523020 474758 523144 474858
rect 523244 474758 523368 474858
rect 523468 474758 523592 474858
rect 523692 474758 523816 474858
rect 523916 474758 523940 474858
rect 517280 474634 523940 474758
rect 517280 474534 517320 474634
rect 517420 474534 517544 474634
rect 517644 474534 517768 474634
rect 517868 474534 517992 474634
rect 518092 474534 518216 474634
rect 518316 474534 518440 474634
rect 518540 474534 518664 474634
rect 518764 474534 518888 474634
rect 518988 474534 519112 474634
rect 519212 474534 519336 474634
rect 519436 474534 519560 474634
rect 519660 474534 519784 474634
rect 519884 474534 520008 474634
rect 520108 474534 520232 474634
rect 520332 474534 520456 474634
rect 520556 474534 520680 474634
rect 520780 474534 520904 474634
rect 521004 474534 521128 474634
rect 521228 474534 521352 474634
rect 521452 474534 521576 474634
rect 521676 474534 521800 474634
rect 521900 474534 522024 474634
rect 522124 474534 522248 474634
rect 522348 474534 522472 474634
rect 522572 474534 522696 474634
rect 522796 474534 522920 474634
rect 523020 474534 523144 474634
rect 523244 474534 523368 474634
rect 523468 474534 523592 474634
rect 523692 474534 523816 474634
rect 523916 474534 523940 474634
rect 517280 474410 523940 474534
rect 517280 474310 517320 474410
rect 517420 474310 517544 474410
rect 517644 474310 517768 474410
rect 517868 474310 517992 474410
rect 518092 474310 518216 474410
rect 518316 474310 518440 474410
rect 518540 474310 518664 474410
rect 518764 474310 518888 474410
rect 518988 474310 519112 474410
rect 519212 474310 519336 474410
rect 519436 474310 519560 474410
rect 519660 474310 519784 474410
rect 519884 474310 520008 474410
rect 520108 474310 520232 474410
rect 520332 474310 520456 474410
rect 520556 474310 520680 474410
rect 520780 474310 520904 474410
rect 521004 474310 521128 474410
rect 521228 474310 521352 474410
rect 521452 474310 521576 474410
rect 521676 474310 521800 474410
rect 521900 474310 522024 474410
rect 522124 474310 522248 474410
rect 522348 474310 522472 474410
rect 522572 474310 522696 474410
rect 522796 474310 522920 474410
rect 523020 474310 523144 474410
rect 523244 474310 523368 474410
rect 523468 474310 523592 474410
rect 523692 474310 523816 474410
rect 523916 474310 523940 474410
rect 517280 474276 523940 474310
rect 527584 474280 528644 474320
rect 500364 474056 501424 474180
rect 500364 473956 500398 474056
rect 500498 473956 500622 474056
rect 500722 473956 500846 474056
rect 500946 473956 501070 474056
rect 501170 473956 501294 474056
rect 501394 473956 501424 474056
rect 500364 473832 501424 473956
rect 500364 473732 500398 473832
rect 500498 473732 500622 473832
rect 500722 473732 500846 473832
rect 500946 473732 501070 473832
rect 501170 473732 501294 473832
rect 501394 473732 501424 473832
rect 500364 473608 501424 473732
rect 500364 473508 500398 473608
rect 500498 473508 500622 473608
rect 500722 473508 500846 473608
rect 500946 473508 501070 473608
rect 501170 473508 501294 473608
rect 501394 473508 501424 473608
rect 500364 473384 501424 473508
rect 500364 473284 500398 473384
rect 500498 473284 500622 473384
rect 500722 473284 500846 473384
rect 500946 473284 501070 473384
rect 501170 473284 501294 473384
rect 501394 473284 501424 473384
rect 500364 473160 501424 473284
rect 500364 473060 500398 473160
rect 500498 473060 500622 473160
rect 500722 473060 500846 473160
rect 500946 473060 501070 473160
rect 501170 473060 501294 473160
rect 501394 473060 501424 473160
rect 500364 472936 501424 473060
rect 500364 472836 500398 472936
rect 500498 472836 500622 472936
rect 500722 472836 500846 472936
rect 500946 472836 501070 472936
rect 501170 472836 501294 472936
rect 501394 472836 501424 472936
rect 500364 472712 501424 472836
rect 500364 472612 500398 472712
rect 500498 472612 500622 472712
rect 500722 472612 500846 472712
rect 500946 472612 501070 472712
rect 501170 472612 501294 472712
rect 501394 472612 501424 472712
rect 500364 472488 501424 472612
rect 527584 474180 527618 474280
rect 527718 474180 527842 474280
rect 527942 474180 528066 474280
rect 528166 474180 528290 474280
rect 528390 474180 528514 474280
rect 528614 474180 528644 474280
rect 527584 474056 528644 474180
rect 527584 473956 527618 474056
rect 527718 473956 527842 474056
rect 527942 473956 528066 474056
rect 528166 473956 528290 474056
rect 528390 473956 528514 474056
rect 528614 473956 528644 474056
rect 527584 473832 528644 473956
rect 527584 473732 527618 473832
rect 527718 473732 527842 473832
rect 527942 473732 528066 473832
rect 528166 473732 528290 473832
rect 528390 473732 528514 473832
rect 528614 473732 528644 473832
rect 527584 473608 528644 473732
rect 527584 473508 527618 473608
rect 527718 473508 527842 473608
rect 527942 473508 528066 473608
rect 528166 473508 528290 473608
rect 528390 473508 528514 473608
rect 528614 473508 528644 473608
rect 527584 473384 528644 473508
rect 527584 473284 527618 473384
rect 527718 473284 527842 473384
rect 527942 473284 528066 473384
rect 528166 473284 528290 473384
rect 528390 473284 528514 473384
rect 528614 473284 528644 473384
rect 527584 473160 528644 473284
rect 527584 473060 527618 473160
rect 527718 473060 527842 473160
rect 527942 473060 528066 473160
rect 528166 473060 528290 473160
rect 528390 473060 528514 473160
rect 528614 473060 528644 473160
rect 527584 472936 528644 473060
rect 527584 472836 527618 472936
rect 527718 472836 527842 472936
rect 527942 472836 528066 472936
rect 528166 472836 528290 472936
rect 528390 472836 528514 472936
rect 528614 472836 528644 472936
rect 527584 472712 528644 472836
rect 527584 472612 527618 472712
rect 527718 472612 527842 472712
rect 527942 472612 528066 472712
rect 528166 472612 528290 472712
rect 528390 472612 528514 472712
rect 528614 472612 528644 472712
rect 500364 472388 500398 472488
rect 500498 472388 500622 472488
rect 500722 472388 500846 472488
rect 500946 472388 501070 472488
rect 501170 472388 501294 472488
rect 501394 472388 501424 472488
rect 500364 472264 501424 472388
rect 525651 472504 526507 472513
rect 506364 472316 506434 472322
rect 500364 472164 500398 472264
rect 500498 472164 500622 472264
rect 500722 472164 500846 472264
rect 500946 472164 501070 472264
rect 501170 472164 501294 472264
rect 501394 472164 501424 472264
rect 500364 472040 501424 472164
rect 500364 471940 500398 472040
rect 500498 471940 500622 472040
rect 500722 471940 500846 472040
rect 500946 471940 501070 472040
rect 501170 471940 501294 472040
rect 501394 471940 501424 472040
rect 500364 471816 501424 471940
rect 500364 471716 500398 471816
rect 500498 471716 500622 471816
rect 500722 471716 500846 471816
rect 500946 471716 501070 471816
rect 501170 471716 501294 471816
rect 501394 471716 501424 471816
rect 500364 471592 501424 471716
rect 500364 471492 500398 471592
rect 500498 471492 500622 471592
rect 500722 471492 500846 471592
rect 500946 471492 501070 471592
rect 501170 471492 501294 471592
rect 501394 471492 501424 471592
rect 500364 471368 501424 471492
rect 500364 471268 500398 471368
rect 500498 471268 500622 471368
rect 500722 471268 500846 471368
rect 500946 471268 501070 471368
rect 501170 471268 501294 471368
rect 501394 471268 501424 471368
rect 500364 471144 501424 471268
rect 500364 471044 500398 471144
rect 500498 471044 500622 471144
rect 500722 471044 500846 471144
rect 500946 471044 501070 471144
rect 501170 471044 501294 471144
rect 501394 471044 501424 471144
rect 500364 470920 501424 471044
rect 500364 470820 500398 470920
rect 500498 470820 500622 470920
rect 500722 470820 500846 470920
rect 500946 470820 501070 470920
rect 501170 470820 501294 470920
rect 501394 470820 501424 470920
rect 500364 470696 501424 470820
rect 500364 470596 500398 470696
rect 500498 470596 500622 470696
rect 500722 470596 500846 470696
rect 500946 470596 501070 470696
rect 501170 470596 501294 470696
rect 501394 470596 501424 470696
rect 500364 470472 501424 470596
rect 500364 470372 500398 470472
rect 500498 470372 500622 470472
rect 500722 470372 500846 470472
rect 500946 470372 501070 470472
rect 501170 470372 501294 470472
rect 501394 470372 501424 470472
rect 500364 470248 501424 470372
rect 500364 470148 500398 470248
rect 500498 470148 500622 470248
rect 500722 470148 500846 470248
rect 500946 470148 501070 470248
rect 501170 470148 501294 470248
rect 501394 470148 501424 470248
rect 506090 471398 506224 472269
rect 506090 471346 506164 471398
rect 506216 471346 506224 471398
rect 500364 470024 501424 470148
rect 500364 469924 500398 470024
rect 500498 469924 500622 470024
rect 500722 469924 500846 470024
rect 500946 469924 501070 470024
rect 501170 469924 501294 470024
rect 501394 469924 501424 470024
rect 500364 469800 501424 469924
rect 502864 470210 502988 470220
rect 500364 469700 500398 469800
rect 500498 469700 500622 469800
rect 500722 469700 500846 469800
rect 500946 469700 501070 469800
rect 501170 469700 501294 469800
rect 501394 469700 501424 469800
rect 500364 469576 501424 469700
rect 500364 469476 500398 469576
rect 500498 469476 500622 469576
rect 500722 469476 500846 469576
rect 500946 469476 501070 469576
rect 501170 469476 501294 469576
rect 501394 469476 501424 469576
rect 500364 469352 501424 469476
rect 500364 469252 500398 469352
rect 500498 469252 500622 469352
rect 500722 469252 500846 469352
rect 500946 469252 501070 469352
rect 501170 469252 501294 469352
rect 501394 469252 501424 469352
rect 500364 469128 501424 469252
rect 500364 469028 500398 469128
rect 500498 469028 500622 469128
rect 500722 469028 500846 469128
rect 500946 469028 501070 469128
rect 501170 469028 501294 469128
rect 501394 469028 501424 469128
rect 500364 468904 501424 469028
rect 500364 468804 500398 468904
rect 500498 468804 500622 468904
rect 500722 468804 500846 468904
rect 500946 468804 501070 468904
rect 501170 468804 501294 468904
rect 501394 468804 501424 468904
rect 500364 468680 501424 468804
rect 500364 468580 500398 468680
rect 500498 468580 500622 468680
rect 500722 468580 500846 468680
rect 500946 468580 501070 468680
rect 501170 468580 501294 468680
rect 501394 468580 501424 468680
rect 500364 468456 501424 468580
rect 500364 468356 500398 468456
rect 500498 468356 500622 468456
rect 500722 468356 500846 468456
rect 500946 468356 501070 468456
rect 501170 468356 501294 468456
rect 501394 468356 501424 468456
rect 500364 468232 501424 468356
rect 500364 468132 500398 468232
rect 500498 468132 500622 468232
rect 500722 468132 500846 468232
rect 500946 468132 501070 468232
rect 501170 468132 501294 468232
rect 501394 468132 501424 468232
rect 500364 468008 501424 468132
rect 500364 467908 500398 468008
rect 500498 467908 500622 468008
rect 500722 467908 500846 468008
rect 500946 467908 501070 468008
rect 501170 467908 501294 468008
rect 501394 467908 501424 468008
rect 500364 467784 501424 467908
rect 500364 467684 500398 467784
rect 500498 467684 500622 467784
rect 500722 467684 500846 467784
rect 500946 467684 501070 467784
rect 501170 467684 501294 467784
rect 501394 467684 501424 467784
rect 500364 467660 501424 467684
rect 502664 469876 502790 469882
rect 502664 469682 502670 469876
rect 502784 469682 502790 469876
rect 502664 469676 502790 469682
rect 502664 468996 502788 469676
rect 502664 468944 502674 468996
rect 502778 468944 502788 468996
rect 502664 468424 502788 468944
rect 502664 468372 502674 468424
rect 502778 468372 502788 468424
rect 502664 467852 502788 468372
rect 502664 467800 502674 467852
rect 502778 467800 502788 467852
rect 500364 463810 501424 463850
rect 500364 463710 500398 463810
rect 500498 463710 500622 463810
rect 500722 463710 500846 463810
rect 500946 463710 501070 463810
rect 501170 463710 501294 463810
rect 501394 463710 501424 463810
rect 500364 463586 501424 463710
rect 500364 463486 500398 463586
rect 500498 463486 500622 463586
rect 500722 463486 500846 463586
rect 500946 463486 501070 463586
rect 501170 463486 501294 463586
rect 501394 463486 501424 463586
rect 500364 463362 501424 463486
rect 500364 463262 500398 463362
rect 500498 463262 500622 463362
rect 500722 463262 500846 463362
rect 500946 463262 501070 463362
rect 501170 463262 501294 463362
rect 501394 463262 501424 463362
rect 500364 463138 501424 463262
rect 500364 463038 500398 463138
rect 500498 463038 500622 463138
rect 500722 463038 500846 463138
rect 500946 463038 501070 463138
rect 501170 463038 501294 463138
rect 501394 463038 501424 463138
rect 500364 462914 501424 463038
rect 500364 462814 500398 462914
rect 500498 462814 500622 462914
rect 500722 462814 500846 462914
rect 500946 462814 501070 462914
rect 501170 462814 501294 462914
rect 501394 462814 501424 462914
rect 500364 462690 501424 462814
rect 500364 462590 500398 462690
rect 500498 462590 500622 462690
rect 500722 462590 500846 462690
rect 500946 462590 501070 462690
rect 501170 462590 501294 462690
rect 501394 462590 501424 462690
rect 502664 463848 502788 467800
rect 502664 463796 502674 463848
rect 502778 463796 502788 463848
rect 502664 463276 502788 463796
rect 502664 463224 502674 463276
rect 502778 463224 502788 463276
rect 502664 462704 502788 463224
rect 502664 462652 502674 462704
rect 502778 462652 502788 462704
rect 502664 462642 502788 462652
rect 500364 462466 501424 462590
rect 500364 462366 500398 462466
rect 500498 462366 500622 462466
rect 500722 462366 500846 462466
rect 500946 462366 501070 462466
rect 501170 462366 501294 462466
rect 501394 462366 501424 462466
rect 500364 462242 501424 462366
rect 500364 462142 500398 462242
rect 500498 462142 500622 462242
rect 500722 462142 500846 462242
rect 500946 462142 501070 462242
rect 501170 462142 501294 462242
rect 501394 462142 501424 462242
rect 500364 462018 501424 462142
rect 500364 461918 500398 462018
rect 500498 461918 500622 462018
rect 500722 461918 500846 462018
rect 500946 461918 501070 462018
rect 501170 461918 501294 462018
rect 501394 461918 501424 462018
rect 500364 461794 501424 461918
rect 500364 461694 500398 461794
rect 500498 461694 500622 461794
rect 500722 461694 500846 461794
rect 500946 461694 501070 461794
rect 501170 461694 501294 461794
rect 501394 461694 501424 461794
rect 500364 461570 501424 461694
rect 500364 461470 500398 461570
rect 500498 461470 500622 461570
rect 500722 461470 500846 461570
rect 500946 461470 501070 461570
rect 501170 461470 501294 461570
rect 501394 461470 501424 461570
rect 500364 461346 501424 461470
rect 500364 461246 500398 461346
rect 500498 461246 500622 461346
rect 500722 461246 500846 461346
rect 500946 461246 501070 461346
rect 501170 461246 501294 461346
rect 501394 461246 501424 461346
rect 500364 461122 501424 461246
rect 500364 461022 500398 461122
rect 500498 461022 500622 461122
rect 500722 461022 500846 461122
rect 500946 461022 501070 461122
rect 501170 461022 501294 461122
rect 501394 461022 501424 461122
rect 500364 460898 501424 461022
rect 502864 460964 502868 470210
rect 502982 460964 502988 470210
rect 505796 469552 506062 469572
rect 505796 468952 505803 469552
rect 506055 468952 506062 469552
rect 505796 468720 506062 468952
rect 505796 468668 505802 468720
rect 506056 468668 506062 468720
rect 505796 468160 506062 468668
rect 505796 468108 505802 468160
rect 506056 468108 506062 468160
rect 505796 467600 506062 468108
rect 505796 467548 505802 467600
rect 506056 467548 506062 467600
rect 505698 467122 505768 467128
rect 505698 466914 505708 467122
rect 505766 466914 505768 467122
rect 505698 466550 505768 466914
rect 505698 466342 505704 466550
rect 505762 466342 505768 466550
rect 505698 466082 505768 466342
rect 505702 465978 505768 466082
rect 505702 465770 505708 465978
rect 505766 465770 505768 465978
rect 505702 465406 505768 465770
rect 505702 465198 505708 465406
rect 505766 465198 505768 465406
rect 505702 464834 505768 465198
rect 505702 464626 505708 464834
rect 505766 464626 505768 464834
rect 505702 464262 505768 464626
rect 505702 464054 505708 464262
rect 505766 464054 505768 464262
rect 505702 464048 505768 464054
rect 505796 466700 506062 467548
rect 505796 466648 505802 466700
rect 506056 466648 506062 466700
rect 505796 465556 506062 466648
rect 505796 465504 505802 465556
rect 506056 465504 506062 465556
rect 505796 464412 506062 465504
rect 505796 464360 505802 464412
rect 506056 464360 506062 464412
rect 502864 460954 502988 460964
rect 505796 463612 506062 464360
rect 506090 466820 506224 471346
rect 506364 472264 506370 472316
rect 506422 472264 506434 472316
rect 506364 470482 506434 472264
rect 506364 470430 506376 470482
rect 506428 470430 506434 470482
rect 506364 469876 506434 470430
rect 506364 469682 506370 469876
rect 506428 469682 506434 469876
rect 506364 469676 506434 469682
rect 509930 470184 512010 470196
rect 509930 470124 509940 470184
rect 510010 470124 510034 470184
rect 510104 470176 512010 470184
rect 510104 470124 511770 470176
rect 509930 470116 511770 470124
rect 511830 470116 511890 470176
rect 511950 470116 512010 470176
rect 509930 470112 512010 470116
rect 509930 470052 509940 470112
rect 510010 470052 510034 470112
rect 510104 470056 512010 470112
rect 510104 470052 511770 470056
rect 509930 470040 511770 470052
rect 509930 469980 509940 470040
rect 510010 469980 510034 470040
rect 510104 469996 511770 470040
rect 511830 469996 511890 470056
rect 511950 469996 512010 470056
rect 510104 469980 512010 469996
rect 509930 469968 512010 469980
rect 509930 469908 509940 469968
rect 510010 469908 510034 469968
rect 510104 469936 512010 469968
rect 510104 469908 511770 469936
rect 509930 469896 511770 469908
rect 509930 469836 509940 469896
rect 510010 469836 510034 469896
rect 510104 469876 511770 469896
rect 511830 469876 511890 469936
rect 511950 469876 512010 469936
rect 510104 469836 512010 469876
rect 509930 469824 512010 469836
rect 509930 469764 509940 469824
rect 510010 469764 510034 469824
rect 510104 469816 512010 469824
rect 510104 469764 511770 469816
rect 509930 469756 511770 469764
rect 511830 469756 511890 469816
rect 511950 469756 512010 469816
rect 509930 469752 512010 469756
rect 509930 469692 509940 469752
rect 510010 469692 510034 469752
rect 510104 469696 512010 469752
rect 510104 469692 511770 469696
rect 509930 469680 511770 469692
rect 509930 469620 509940 469680
rect 510010 469620 510034 469680
rect 510104 469636 511770 469680
rect 511830 469636 511890 469696
rect 511950 469636 512010 469696
rect 510104 469620 512010 469636
rect 509930 469606 512010 469620
rect 506090 466768 506102 466820
rect 506206 466768 506224 466820
rect 506090 466248 506224 466768
rect 506090 466196 506102 466248
rect 506206 466196 506224 466248
rect 506090 465676 506224 466196
rect 506090 465624 506102 465676
rect 506206 465624 506224 465676
rect 506090 465104 506224 465624
rect 506090 465052 506102 465104
rect 506206 465052 506224 465104
rect 506090 464532 506224 465052
rect 506090 464480 506102 464532
rect 506206 464480 506224 464532
rect 506090 463960 506224 464480
rect 506090 463908 506102 463960
rect 506206 463908 506224 463960
rect 506090 463898 506224 463908
rect 508212 467088 508292 467108
rect 508212 466944 508218 467088
rect 508272 466944 508292 467088
rect 508212 465944 508292 466944
rect 508212 465800 508218 465944
rect 508272 465800 508292 465944
rect 508212 464800 508292 465800
rect 508212 464656 508218 464800
rect 508272 464656 508292 464800
rect 505796 463560 505802 463612
rect 506056 463560 506062 463612
rect 505796 463052 506062 463560
rect 505796 463000 505802 463052
rect 506056 463000 506062 463052
rect 505796 462492 506062 463000
rect 505796 462440 505802 462492
rect 506056 462440 506062 462492
rect 505796 461061 506062 462440
rect 508212 461310 508292 464656
rect 508212 461194 508292 461200
rect 508352 466516 508432 466536
rect 508352 466372 508358 466516
rect 508412 466372 508432 466516
rect 508352 465372 508432 466372
rect 508352 465228 508358 465372
rect 508412 465228 508432 465372
rect 508352 464228 508432 465228
rect 508352 464084 508358 464228
rect 508412 464084 508432 464228
rect 500364 460798 500398 460898
rect 500498 460798 500622 460898
rect 500722 460798 500846 460898
rect 500946 460798 501070 460898
rect 501170 460798 501294 460898
rect 501394 460798 501424 460898
rect 500364 460674 501424 460798
rect 500364 460574 500398 460674
rect 500498 460574 500622 460674
rect 500722 460574 500846 460674
rect 500946 460574 501070 460674
rect 501170 460574 501294 460674
rect 501394 460574 501424 460674
rect 500364 460450 501424 460574
rect 505796 460461 505803 461061
rect 506055 460461 506062 461061
rect 508352 460854 508432 464084
rect 508352 460728 508432 460734
rect 511228 461310 511828 461316
rect 511228 461190 511532 461310
rect 511824 461190 511828 461310
rect 525651 461248 525660 472504
rect 526498 461248 526507 472504
rect 527584 472488 528644 472612
rect 527584 472388 527618 472488
rect 527718 472388 527842 472488
rect 527942 472388 528066 472488
rect 528166 472388 528290 472488
rect 528390 472388 528514 472488
rect 528614 472388 528644 472488
rect 527584 472264 528644 472388
rect 527584 472164 527618 472264
rect 527718 472164 527842 472264
rect 527942 472164 528066 472264
rect 528166 472164 528290 472264
rect 528390 472164 528514 472264
rect 528614 472164 528644 472264
rect 527584 472040 528644 472164
rect 527584 471940 527618 472040
rect 527718 471940 527842 472040
rect 527942 471940 528066 472040
rect 528166 471940 528290 472040
rect 528390 471940 528514 472040
rect 528614 471940 528644 472040
rect 527584 471816 528644 471940
rect 527584 471716 527618 471816
rect 527718 471716 527842 471816
rect 527942 471716 528066 471816
rect 528166 471716 528290 471816
rect 528390 471716 528514 471816
rect 528614 471716 528644 471816
rect 527584 471592 528644 471716
rect 527584 471492 527618 471592
rect 527718 471492 527842 471592
rect 527942 471492 528066 471592
rect 528166 471492 528290 471592
rect 528390 471492 528514 471592
rect 528614 471492 528644 471592
rect 527584 471368 528644 471492
rect 527584 471268 527618 471368
rect 527718 471268 527842 471368
rect 527942 471268 528066 471368
rect 528166 471268 528290 471368
rect 528390 471268 528514 471368
rect 528614 471268 528644 471368
rect 527584 471144 528644 471268
rect 527584 471044 527618 471144
rect 527718 471044 527842 471144
rect 527942 471044 528066 471144
rect 528166 471044 528290 471144
rect 528390 471044 528514 471144
rect 528614 471044 528644 471144
rect 527584 470920 528644 471044
rect 527584 470820 527618 470920
rect 527718 470820 527842 470920
rect 527942 470820 528066 470920
rect 528166 470820 528290 470920
rect 528390 470820 528514 470920
rect 528614 470820 528644 470920
rect 527584 470696 528644 470820
rect 527584 470596 527618 470696
rect 527718 470596 527842 470696
rect 527942 470596 528066 470696
rect 528166 470596 528290 470696
rect 528390 470596 528514 470696
rect 528614 470596 528644 470696
rect 527584 470472 528644 470596
rect 527584 470372 527618 470472
rect 527718 470372 527842 470472
rect 527942 470372 528066 470472
rect 528166 470372 528290 470472
rect 528390 470372 528514 470472
rect 528614 470372 528644 470472
rect 527584 470248 528644 470372
rect 527584 470148 527618 470248
rect 527718 470148 527842 470248
rect 527942 470148 528066 470248
rect 528166 470148 528290 470248
rect 528390 470148 528514 470248
rect 528614 470148 528644 470248
rect 527584 470024 528644 470148
rect 527584 469924 527618 470024
rect 527718 469924 527842 470024
rect 527942 469924 528066 470024
rect 528166 469924 528290 470024
rect 528390 469924 528514 470024
rect 528614 469924 528644 470024
rect 527584 469800 528644 469924
rect 527584 469700 527618 469800
rect 527718 469700 527842 469800
rect 527942 469700 528066 469800
rect 528166 469700 528290 469800
rect 528390 469700 528514 469800
rect 528614 469700 528644 469800
rect 527584 469576 528644 469700
rect 527584 469476 527618 469576
rect 527718 469476 527842 469576
rect 527942 469476 528066 469576
rect 528166 469476 528290 469576
rect 528390 469476 528514 469576
rect 528614 469476 528644 469576
rect 527584 469352 528644 469476
rect 527584 469252 527618 469352
rect 527718 469252 527842 469352
rect 527942 469252 528066 469352
rect 528166 469252 528290 469352
rect 528390 469252 528514 469352
rect 528614 469252 528644 469352
rect 527584 469128 528644 469252
rect 527584 469028 527618 469128
rect 527718 469028 527842 469128
rect 527942 469028 528066 469128
rect 528166 469028 528290 469128
rect 528390 469028 528514 469128
rect 528614 469028 528644 469128
rect 527584 468904 528644 469028
rect 527584 468804 527618 468904
rect 527718 468804 527842 468904
rect 527942 468804 528066 468904
rect 528166 468804 528290 468904
rect 528390 468804 528514 468904
rect 528614 468804 528644 468904
rect 527584 468680 528644 468804
rect 527584 468580 527618 468680
rect 527718 468580 527842 468680
rect 527942 468580 528066 468680
rect 528166 468580 528290 468680
rect 528390 468580 528514 468680
rect 528614 468580 528644 468680
rect 527584 468456 528644 468580
rect 527584 468356 527618 468456
rect 527718 468356 527842 468456
rect 527942 468356 528066 468456
rect 528166 468356 528290 468456
rect 528390 468356 528514 468456
rect 528614 468356 528644 468456
rect 527584 468232 528644 468356
rect 527584 468132 527618 468232
rect 527718 468132 527842 468232
rect 527942 468132 528066 468232
rect 528166 468132 528290 468232
rect 528390 468132 528514 468232
rect 528614 468132 528644 468232
rect 527584 468008 528644 468132
rect 527584 467908 527618 468008
rect 527718 467908 527842 468008
rect 527942 467908 528066 468008
rect 528166 467908 528290 468008
rect 528390 467908 528514 468008
rect 528614 467908 528644 468008
rect 527584 467784 528644 467908
rect 527584 467684 527618 467784
rect 527718 467684 527842 467784
rect 527942 467684 528066 467784
rect 528166 467684 528290 467784
rect 528390 467684 528514 467784
rect 528614 467684 528644 467784
rect 527584 467660 528644 467684
rect 525651 461239 526507 461248
rect 527584 463810 528644 463850
rect 527584 463710 527618 463810
rect 527718 463710 527842 463810
rect 527942 463710 528066 463810
rect 528166 463710 528290 463810
rect 528390 463710 528514 463810
rect 528614 463710 528644 463810
rect 527584 463586 528644 463710
rect 527584 463486 527618 463586
rect 527718 463486 527842 463586
rect 527942 463486 528066 463586
rect 528166 463486 528290 463586
rect 528390 463486 528514 463586
rect 528614 463486 528644 463586
rect 527584 463362 528644 463486
rect 527584 463262 527618 463362
rect 527718 463262 527842 463362
rect 527942 463262 528066 463362
rect 528166 463262 528290 463362
rect 528390 463262 528514 463362
rect 528614 463262 528644 463362
rect 527584 463138 528644 463262
rect 527584 463038 527618 463138
rect 527718 463038 527842 463138
rect 527942 463038 528066 463138
rect 528166 463038 528290 463138
rect 528390 463038 528514 463138
rect 528614 463038 528644 463138
rect 527584 462914 528644 463038
rect 527584 462814 527618 462914
rect 527718 462814 527842 462914
rect 527942 462814 528066 462914
rect 528166 462814 528290 462914
rect 528390 462814 528514 462914
rect 528614 462814 528644 462914
rect 527584 462690 528644 462814
rect 527584 462590 527618 462690
rect 527718 462590 527842 462690
rect 527942 462590 528066 462690
rect 528166 462590 528290 462690
rect 528390 462590 528514 462690
rect 528614 462590 528644 462690
rect 527584 462466 528644 462590
rect 527584 462366 527618 462466
rect 527718 462366 527842 462466
rect 527942 462366 528066 462466
rect 528166 462366 528290 462466
rect 528390 462366 528514 462466
rect 528614 462366 528644 462466
rect 527584 462242 528644 462366
rect 527584 462142 527618 462242
rect 527718 462142 527842 462242
rect 527942 462142 528066 462242
rect 528166 462142 528290 462242
rect 528390 462142 528514 462242
rect 528614 462142 528644 462242
rect 527584 462018 528644 462142
rect 527584 461918 527618 462018
rect 527718 461918 527842 462018
rect 527942 461918 528066 462018
rect 528166 461918 528290 462018
rect 528390 461918 528514 462018
rect 528614 461918 528644 462018
rect 527584 461794 528644 461918
rect 527584 461694 527618 461794
rect 527718 461694 527842 461794
rect 527942 461694 528066 461794
rect 528166 461694 528290 461794
rect 528390 461694 528514 461794
rect 528614 461694 528644 461794
rect 527584 461570 528644 461694
rect 527584 461470 527618 461570
rect 527718 461470 527842 461570
rect 527942 461470 528066 461570
rect 528166 461470 528290 461570
rect 528390 461470 528514 461570
rect 528614 461470 528644 461570
rect 527584 461346 528644 461470
rect 527584 461246 527618 461346
rect 527718 461246 527842 461346
rect 527942 461246 528066 461346
rect 528166 461246 528290 461346
rect 528390 461246 528514 461346
rect 528614 461246 528644 461346
rect 500364 460350 500398 460450
rect 500498 460350 500622 460450
rect 500722 460350 500846 460450
rect 500946 460350 501070 460450
rect 501170 460350 501294 460450
rect 501394 460350 501424 460450
rect 500364 460226 501424 460350
rect 500364 460126 500398 460226
rect 500498 460126 500622 460226
rect 500722 460126 500846 460226
rect 500946 460126 501070 460226
rect 501170 460126 501294 460226
rect 501394 460126 501424 460226
rect 500364 460002 501424 460126
rect 500364 459902 500398 460002
rect 500498 459902 500622 460002
rect 500722 459902 500846 460002
rect 500946 459902 501070 460002
rect 501170 459902 501294 460002
rect 501394 459902 501424 460002
rect 500364 459778 501424 459902
rect 500364 459678 500398 459778
rect 500498 459678 500622 459778
rect 500722 459678 500846 459778
rect 500946 459678 501070 459778
rect 501170 459678 501294 459778
rect 501394 459678 501424 459778
rect 500364 459554 501424 459678
rect 500364 459454 500398 459554
rect 500498 459454 500622 459554
rect 500722 459454 500846 459554
rect 500946 459454 501070 459554
rect 501170 459454 501294 459554
rect 501394 459454 501424 459554
rect 500364 459330 501424 459454
rect 500364 459230 500398 459330
rect 500498 459230 500622 459330
rect 500722 459230 500846 459330
rect 500946 459230 501070 459330
rect 501170 459230 501294 459330
rect 501394 459230 501424 459330
rect 500364 459106 501424 459230
rect 500364 459006 500398 459106
rect 500498 459006 500622 459106
rect 500722 459006 500846 459106
rect 500946 459006 501070 459106
rect 501170 459006 501294 459106
rect 501394 459006 501424 459106
rect 500364 458882 501424 459006
rect 500364 458782 500398 458882
rect 500498 458782 500622 458882
rect 500722 458782 500846 458882
rect 500946 458782 501070 458882
rect 501170 458782 501294 458882
rect 501394 458782 501424 458882
rect 500364 458658 501424 458782
rect 500364 458558 500398 458658
rect 500498 458558 500622 458658
rect 500722 458558 500846 458658
rect 500946 458558 501070 458658
rect 501170 458558 501294 458658
rect 501394 458558 501424 458658
rect 500364 458434 501424 458558
rect 500364 458334 500398 458434
rect 500498 458334 500622 458434
rect 500722 458334 500846 458434
rect 500946 458334 501070 458434
rect 501170 458334 501294 458434
rect 501394 458334 501424 458434
rect 500364 458210 501424 458334
rect 500364 458110 500398 458210
rect 500498 458110 500622 458210
rect 500722 458110 500846 458210
rect 500946 458110 501070 458210
rect 501170 458110 501294 458210
rect 501394 458110 501424 458210
rect 500364 457986 501424 458110
rect 500364 457886 500398 457986
rect 500498 457886 500622 457986
rect 500722 457886 500846 457986
rect 500946 457886 501070 457986
rect 501170 457886 501294 457986
rect 501394 457886 501424 457986
rect 500364 457762 501424 457886
rect 500364 457662 500398 457762
rect 500498 457662 500622 457762
rect 500722 457662 500846 457762
rect 500946 457662 501070 457762
rect 501170 457662 501294 457762
rect 501394 457662 501424 457762
rect 500364 457538 501424 457662
rect 500364 457438 500398 457538
rect 500498 457438 500622 457538
rect 500722 457438 500846 457538
rect 500946 457438 501070 457538
rect 501170 457438 501294 457538
rect 501394 457438 501424 457538
rect 500364 457314 501424 457438
rect 500364 457214 500398 457314
rect 500498 457214 500622 457314
rect 500722 457214 500846 457314
rect 500946 457214 501070 457314
rect 501170 457214 501294 457314
rect 501394 457214 501424 457314
rect 500364 457190 501424 457214
rect 502424 460446 502760 460456
rect 502424 442508 502432 460446
rect 502750 458882 502760 460446
rect 502808 460442 502968 460448
rect 502808 459974 502814 460442
rect 502962 459974 502968 460442
rect 502808 459122 502968 459974
rect 505796 460442 506062 460461
rect 505796 459974 505802 460442
rect 506056 459974 506062 460442
rect 505796 459968 506062 459974
rect 502808 458982 502828 459122
rect 502948 458982 502968 459122
rect 502750 458762 502768 458882
rect 502750 457962 502760 458762
rect 502808 458662 502968 458982
rect 502808 458522 502828 458662
rect 502948 458522 502968 458662
rect 502808 458202 502968 458522
rect 502808 458062 502828 458202
rect 502948 458062 502968 458202
rect 502750 457842 502768 457962
rect 502750 457042 502760 457842
rect 502808 457742 502968 458062
rect 502808 457602 502828 457742
rect 502948 457602 502968 457742
rect 502808 457282 502968 457602
rect 502808 457142 502828 457282
rect 502948 457142 502968 457282
rect 502750 456922 502768 457042
rect 502750 456122 502760 456922
rect 502808 456822 502968 457142
rect 502808 456682 502828 456822
rect 502948 456682 502968 456822
rect 502808 456362 502968 456682
rect 502808 456222 502828 456362
rect 502948 456222 502968 456362
rect 502750 456002 502768 456122
rect 502750 455202 502760 456002
rect 502808 455902 502968 456222
rect 502808 455762 502828 455902
rect 502948 455762 502968 455902
rect 502808 455442 502968 455762
rect 502808 455302 502828 455442
rect 502948 455302 502968 455442
rect 502750 455082 502768 455202
rect 502750 453382 502760 455082
rect 502808 454982 502968 455302
rect 502808 454842 502828 454982
rect 502948 454842 502968 454982
rect 502808 453622 502968 454842
rect 502808 453482 502828 453622
rect 502948 453482 502968 453622
rect 502750 453262 502768 453382
rect 502750 452462 502760 453262
rect 502808 453162 502968 453482
rect 502808 453022 502828 453162
rect 502948 453022 502968 453162
rect 502808 452702 502968 453022
rect 502808 452562 502828 452702
rect 502948 452562 502968 452702
rect 502750 452342 502768 452462
rect 502750 451542 502760 452342
rect 502808 452242 502968 452562
rect 502808 452102 502828 452242
rect 502948 452102 502968 452242
rect 502808 451782 502968 452102
rect 502808 451642 502828 451782
rect 502948 451642 502968 451782
rect 502750 451422 502768 451542
rect 502750 450622 502760 451422
rect 502808 451322 502968 451642
rect 502808 451182 502828 451322
rect 502948 451182 502968 451322
rect 502808 450862 502968 451182
rect 502808 450722 502828 450862
rect 502948 450722 502968 450862
rect 502750 450502 502768 450622
rect 502750 449702 502760 450502
rect 502808 450402 502968 450722
rect 502808 450262 502828 450402
rect 502948 450262 502968 450402
rect 502808 449942 502968 450262
rect 502808 449802 502828 449942
rect 502948 449802 502968 449942
rect 502750 449582 502768 449702
rect 502750 447882 502760 449582
rect 502808 449482 502968 449802
rect 502808 449342 502828 449482
rect 502948 449342 502968 449482
rect 502808 448122 502968 449342
rect 502808 447982 502828 448122
rect 502948 447982 502968 448122
rect 502750 447762 502768 447882
rect 502750 446962 502760 447762
rect 502808 447662 502968 447982
rect 502808 447522 502828 447662
rect 502948 447522 502968 447662
rect 502808 447202 502968 447522
rect 502808 447062 502828 447202
rect 502948 447062 502968 447202
rect 502750 446842 502768 446962
rect 502750 446042 502760 446842
rect 502808 446742 502968 447062
rect 502808 446602 502828 446742
rect 502948 446602 502968 446742
rect 502808 446282 502968 446602
rect 502808 446142 502828 446282
rect 502948 446142 502968 446282
rect 502750 445922 502768 446042
rect 502750 445122 502760 445922
rect 502808 445822 502968 446142
rect 502808 445682 502828 445822
rect 502948 445682 502968 445822
rect 502808 445362 502968 445682
rect 502808 445222 502828 445362
rect 502948 445222 502968 445362
rect 502750 445002 502768 445122
rect 502750 444202 502760 445002
rect 502808 444902 502968 445222
rect 502808 444762 502828 444902
rect 502948 444762 502968 444902
rect 502808 444442 502968 444762
rect 502808 444302 502828 444442
rect 502948 444302 502968 444442
rect 502750 444082 502768 444202
rect 502750 442508 502760 444082
rect 502808 443982 502968 444302
rect 502808 443842 502828 443982
rect 502948 443842 502968 443982
rect 502808 443822 502968 443842
rect 511228 456636 511828 461190
rect 527584 461122 528644 461246
rect 527584 461022 527618 461122
rect 527718 461022 527842 461122
rect 527942 461022 528066 461122
rect 528166 461022 528290 461122
rect 528390 461022 528514 461122
rect 528614 461022 528644 461122
rect 527584 460898 528644 461022
rect 512110 460858 512536 460860
rect 512110 460854 513294 460858
rect 512110 460734 512116 460854
rect 512530 460734 513294 460854
rect 512110 460728 513294 460734
rect 511228 454648 511534 456636
rect 511822 454648 511828 456636
rect 511228 448336 511828 454648
rect 511228 446348 511534 448336
rect 511822 446348 511828 448336
rect 502424 442498 502760 442508
rect 502426 442486 502726 442498
rect 503646 441668 504594 441674
rect 503646 440732 503652 441668
rect 504588 440732 504594 441668
rect 500384 437540 501444 437580
rect 500384 437440 500418 437540
rect 500518 437440 500642 437540
rect 500742 437440 500866 437540
rect 500966 437440 501090 437540
rect 501190 437440 501314 437540
rect 501414 437440 501444 437540
rect 500384 437316 501444 437440
rect 500384 437216 500418 437316
rect 500518 437216 500642 437316
rect 500742 437216 500866 437316
rect 500966 437216 501090 437316
rect 501190 437216 501314 437316
rect 501414 437216 501444 437316
rect 500384 437092 501444 437216
rect 500384 436992 500418 437092
rect 500518 436992 500642 437092
rect 500742 436992 500866 437092
rect 500966 436992 501090 437092
rect 501190 436992 501314 437092
rect 501414 436992 501444 437092
rect 500384 436868 501444 436992
rect 500384 436768 500418 436868
rect 500518 436768 500642 436868
rect 500742 436768 500866 436868
rect 500966 436768 501090 436868
rect 501190 436768 501314 436868
rect 501414 436768 501444 436868
rect 500384 436644 501444 436768
rect 500384 436544 500418 436644
rect 500518 436544 500642 436644
rect 500742 436544 500866 436644
rect 500966 436544 501090 436644
rect 501190 436544 501314 436644
rect 501414 436544 501444 436644
rect 500384 436420 501444 436544
rect 500384 436320 500418 436420
rect 500518 436320 500642 436420
rect 500742 436320 500866 436420
rect 500966 436320 501090 436420
rect 501190 436320 501314 436420
rect 501414 436320 501444 436420
rect 500384 436196 501444 436320
rect 500384 436096 500418 436196
rect 500518 436096 500642 436196
rect 500742 436096 500866 436196
rect 500966 436096 501090 436196
rect 501190 436096 501314 436196
rect 501414 436096 501444 436196
rect 503646 436848 504594 440732
rect 503646 436796 503716 436848
rect 503768 436796 503820 436848
rect 503872 436796 503924 436848
rect 503976 436796 504028 436848
rect 504080 436796 504132 436848
rect 504184 436796 504236 436848
rect 504288 436796 504594 436848
rect 503646 436744 504594 436796
rect 503646 436692 503716 436744
rect 503768 436692 503820 436744
rect 503872 436692 503924 436744
rect 503976 436692 504028 436744
rect 504080 436692 504132 436744
rect 504184 436692 504236 436744
rect 504288 436692 504594 436744
rect 503646 436640 504594 436692
rect 503646 436588 503716 436640
rect 503768 436588 503820 436640
rect 503872 436588 503924 436640
rect 503976 436588 504028 436640
rect 504080 436588 504132 436640
rect 504184 436588 504236 436640
rect 504288 436588 504594 436640
rect 503646 436536 504594 436588
rect 503646 436484 503716 436536
rect 503768 436484 503820 436536
rect 503872 436484 503924 436536
rect 503976 436484 504028 436536
rect 504080 436484 504132 436536
rect 504184 436484 504236 436536
rect 504288 436484 504594 436536
rect 503646 436432 504594 436484
rect 503646 436380 503716 436432
rect 503768 436380 503820 436432
rect 503872 436380 503924 436432
rect 503976 436380 504028 436432
rect 504080 436380 504132 436432
rect 504184 436380 504236 436432
rect 504288 436380 504594 436432
rect 503646 436328 504594 436380
rect 503646 436276 503716 436328
rect 503768 436276 503820 436328
rect 503872 436276 503924 436328
rect 503976 436276 504028 436328
rect 504080 436276 504132 436328
rect 504184 436276 504236 436328
rect 504288 436276 504594 436328
rect 503646 436184 504594 436276
rect 508800 440324 509504 440330
rect 508800 439632 508806 440324
rect 509498 439632 509504 440324
rect 500384 435972 501444 436096
rect 500384 435872 500418 435972
rect 500518 435872 500642 435972
rect 500742 435872 500866 435972
rect 500966 435872 501090 435972
rect 501190 435872 501314 435972
rect 501414 435872 501444 435972
rect 500384 435748 501444 435872
rect 500384 435648 500418 435748
rect 500518 435648 500642 435748
rect 500742 435648 500866 435748
rect 500966 435648 501090 435748
rect 501190 435648 501314 435748
rect 501414 435648 501444 435748
rect 500384 435524 501444 435648
rect 500384 435424 500418 435524
rect 500518 435424 500642 435524
rect 500742 435424 500866 435524
rect 500966 435424 501090 435524
rect 501190 435424 501314 435524
rect 501414 435424 501444 435524
rect 500384 435300 501444 435424
rect 500384 435200 500418 435300
rect 500518 435200 500642 435300
rect 500742 435200 500866 435300
rect 500966 435200 501090 435300
rect 501190 435200 501314 435300
rect 501414 435200 501444 435300
rect 500384 435076 501444 435200
rect 500384 434976 500418 435076
rect 500518 434976 500642 435076
rect 500742 434976 500866 435076
rect 500966 434976 501090 435076
rect 501190 434976 501314 435076
rect 501414 434976 501444 435076
rect 500384 434852 501444 434976
rect 508800 435560 509504 439632
rect 511228 439504 511828 446348
rect 512112 460204 513294 460728
rect 512112 459336 512228 460204
rect 513212 459336 513294 460204
rect 512112 457348 512134 459336
rect 513286 457348 513294 459336
rect 512112 445636 512228 457348
rect 513212 445636 513294 457348
rect 527584 460798 527618 460898
rect 527718 460798 527842 460898
rect 527942 460798 528066 460898
rect 528166 460798 528290 460898
rect 528390 460798 528514 460898
rect 528614 460798 528644 460898
rect 527584 460674 528644 460798
rect 527584 460574 527618 460674
rect 527718 460574 527842 460674
rect 527942 460574 528066 460674
rect 528166 460574 528290 460674
rect 528390 460574 528514 460674
rect 528614 460574 528644 460674
rect 527584 460450 528644 460574
rect 527584 460350 527618 460450
rect 527718 460350 527842 460450
rect 527942 460350 528066 460450
rect 528166 460350 528290 460450
rect 528390 460350 528514 460450
rect 528614 460350 528644 460450
rect 527584 460226 528644 460350
rect 527584 460126 527618 460226
rect 527718 460126 527842 460226
rect 527942 460126 528066 460226
rect 528166 460126 528290 460226
rect 528390 460126 528514 460226
rect 528614 460126 528644 460226
rect 527584 460002 528644 460126
rect 527584 459902 527618 460002
rect 527718 459902 527842 460002
rect 527942 459902 528066 460002
rect 528166 459902 528290 460002
rect 528390 459902 528514 460002
rect 528614 459902 528644 460002
rect 527584 459778 528644 459902
rect 527584 459678 527618 459778
rect 527718 459678 527842 459778
rect 527942 459678 528066 459778
rect 528166 459678 528290 459778
rect 528390 459678 528514 459778
rect 528614 459678 528644 459778
rect 527584 459554 528644 459678
rect 527584 459454 527618 459554
rect 527718 459454 527842 459554
rect 527942 459454 528066 459554
rect 528166 459454 528290 459554
rect 528390 459454 528514 459554
rect 528614 459454 528644 459554
rect 527584 459330 528644 459454
rect 527584 459230 527618 459330
rect 527718 459230 527842 459330
rect 527942 459230 528066 459330
rect 528166 459230 528290 459330
rect 528390 459230 528514 459330
rect 528614 459230 528644 459330
rect 527584 459106 528644 459230
rect 527584 459006 527618 459106
rect 527718 459006 527842 459106
rect 527942 459006 528066 459106
rect 528166 459006 528290 459106
rect 528390 459006 528514 459106
rect 528614 459006 528644 459106
rect 527584 458882 528644 459006
rect 527584 458782 527618 458882
rect 527718 458782 527842 458882
rect 527942 458782 528066 458882
rect 528166 458782 528290 458882
rect 528390 458782 528514 458882
rect 528614 458782 528644 458882
rect 527584 458658 528644 458782
rect 527584 458558 527618 458658
rect 527718 458558 527842 458658
rect 527942 458558 528066 458658
rect 528166 458558 528290 458658
rect 528390 458558 528514 458658
rect 528614 458558 528644 458658
rect 527584 458434 528644 458558
rect 527584 458334 527618 458434
rect 527718 458334 527842 458434
rect 527942 458334 528066 458434
rect 528166 458334 528290 458434
rect 528390 458334 528514 458434
rect 528614 458334 528644 458434
rect 527584 458210 528644 458334
rect 527584 458110 527618 458210
rect 527718 458110 527842 458210
rect 527942 458110 528066 458210
rect 528166 458110 528290 458210
rect 528390 458110 528514 458210
rect 528614 458110 528644 458210
rect 527584 457986 528644 458110
rect 527584 457886 527618 457986
rect 527718 457886 527842 457986
rect 527942 457886 528066 457986
rect 528166 457886 528290 457986
rect 528390 457886 528514 457986
rect 528614 457886 528644 457986
rect 527584 457762 528644 457886
rect 527584 457662 527618 457762
rect 527718 457662 527842 457762
rect 527942 457662 528066 457762
rect 528166 457662 528290 457762
rect 528390 457662 528514 457762
rect 528614 457662 528644 457762
rect 527584 457538 528644 457662
rect 527584 457438 527618 457538
rect 527718 457438 527842 457538
rect 527942 457438 528066 457538
rect 528166 457438 528290 457538
rect 528390 457438 528514 457538
rect 528614 457438 528644 457538
rect 527584 457314 528644 457438
rect 527584 457214 527618 457314
rect 527718 457214 527842 457314
rect 527942 457214 528066 457314
rect 528166 457214 528290 457314
rect 528390 457214 528514 457314
rect 528614 457214 528644 457314
rect 527584 457190 528644 457214
rect 522988 455788 524158 455794
rect 522988 455230 522994 455788
rect 523414 455230 523594 455788
rect 524152 455230 524158 455788
rect 522988 455224 524158 455230
rect 562380 455440 567480 455520
rect 562380 455360 562480 455440
rect 562560 455360 562640 455440
rect 562720 455360 562800 455440
rect 562880 455360 562960 455440
rect 563040 455360 563120 455440
rect 563200 455360 563280 455440
rect 563360 455360 563440 455440
rect 563520 455360 563600 455440
rect 563680 455360 563760 455440
rect 563840 455360 563920 455440
rect 564000 455360 564080 455440
rect 564160 455360 564240 455440
rect 564320 455360 564400 455440
rect 564480 455360 564560 455440
rect 564640 455360 564720 455440
rect 564800 455360 564880 455440
rect 564960 455360 565040 455440
rect 565120 455360 565200 455440
rect 565280 455360 565360 455440
rect 565440 455360 565520 455440
rect 565600 455360 565680 455440
rect 565760 455360 565840 455440
rect 565920 455360 566000 455440
rect 566080 455360 566160 455440
rect 566240 455360 566320 455440
rect 566400 455360 566480 455440
rect 566560 455360 566640 455440
rect 566720 455360 566800 455440
rect 566880 455360 566960 455440
rect 567040 455360 567120 455440
rect 567200 455360 567280 455440
rect 567360 455360 567480 455440
rect 562380 455280 567480 455360
rect 562380 455200 562480 455280
rect 562560 455200 562640 455280
rect 562720 455200 562800 455280
rect 562880 455200 562960 455280
rect 563040 455200 563120 455280
rect 563200 455200 563280 455280
rect 563360 455200 563440 455280
rect 563520 455200 563600 455280
rect 563680 455200 563760 455280
rect 563840 455200 563920 455280
rect 564000 455200 564080 455280
rect 564160 455200 564240 455280
rect 564320 455200 564400 455280
rect 564480 455200 564560 455280
rect 564640 455200 564720 455280
rect 564800 455200 564880 455280
rect 564960 455200 565040 455280
rect 565120 455200 565200 455280
rect 565280 455200 565360 455280
rect 565440 455200 565520 455280
rect 565600 455200 565680 455280
rect 565760 455200 565840 455280
rect 565920 455200 566000 455280
rect 566080 455200 566160 455280
rect 566240 455200 566320 455280
rect 566400 455200 566480 455280
rect 566560 455200 566640 455280
rect 566720 455200 566800 455280
rect 566880 455200 566960 455280
rect 567040 455200 567120 455280
rect 567200 455200 567280 455280
rect 567360 455200 567480 455280
rect 562380 455160 567480 455200
rect 572540 455440 577640 455520
rect 572540 455360 572640 455440
rect 572720 455360 572800 455440
rect 572880 455360 572960 455440
rect 573040 455360 573120 455440
rect 573200 455360 573280 455440
rect 573360 455360 573440 455440
rect 573520 455360 573600 455440
rect 573680 455360 573760 455440
rect 573840 455360 573920 455440
rect 574000 455360 574080 455440
rect 574160 455360 574240 455440
rect 574320 455360 574400 455440
rect 574480 455360 574560 455440
rect 574640 455360 574720 455440
rect 574800 455360 574880 455440
rect 574960 455360 575040 455440
rect 575120 455360 575200 455440
rect 575280 455360 575360 455440
rect 575440 455360 575520 455440
rect 575600 455360 575680 455440
rect 575760 455360 575840 455440
rect 575920 455360 576000 455440
rect 576080 455360 576160 455440
rect 576240 455360 576320 455440
rect 576400 455360 576480 455440
rect 576560 455360 576640 455440
rect 576720 455360 576800 455440
rect 576880 455360 576960 455440
rect 577040 455360 577120 455440
rect 577200 455360 577280 455440
rect 577360 455360 577440 455440
rect 577520 455360 577640 455440
rect 572540 455280 577640 455360
rect 572540 455200 572640 455280
rect 572720 455200 572800 455280
rect 572880 455200 572960 455280
rect 573040 455200 573120 455280
rect 573200 455200 573280 455280
rect 573360 455200 573440 455280
rect 573520 455200 573600 455280
rect 573680 455200 573760 455280
rect 573840 455200 573920 455280
rect 574000 455200 574080 455280
rect 574160 455200 574240 455280
rect 574320 455200 574400 455280
rect 574480 455200 574560 455280
rect 574640 455200 574720 455280
rect 574800 455200 574880 455280
rect 574960 455200 575040 455280
rect 575120 455200 575200 455280
rect 575280 455200 575360 455280
rect 575440 455200 575520 455280
rect 575600 455200 575680 455280
rect 575760 455200 575840 455280
rect 575920 455200 576000 455280
rect 576080 455200 576160 455280
rect 576240 455200 576320 455280
rect 576400 455200 576480 455280
rect 576560 455200 576640 455280
rect 576720 455200 576800 455280
rect 576880 455200 576960 455280
rect 577040 455200 577120 455280
rect 577200 455200 577280 455280
rect 577360 455200 577440 455280
rect 577520 455200 577640 455280
rect 572540 455160 577640 455200
rect 522188 454970 523420 454976
rect 522188 454412 522198 454970
rect 522690 454412 522994 454970
rect 523414 454412 523420 454970
rect 522188 454406 523420 454412
rect 562102 453919 567622 453979
rect 562102 453859 562222 453919
rect 562282 453859 562342 453919
rect 562402 453859 562462 453919
rect 562522 453859 562582 453919
rect 562642 453859 562702 453919
rect 562762 453859 562822 453919
rect 562882 453859 562942 453919
rect 563002 453859 563062 453919
rect 563122 453859 563182 453919
rect 563242 453859 563302 453919
rect 563362 453859 563422 453919
rect 563482 453859 563542 453919
rect 563602 453859 563662 453919
rect 563722 453859 563782 453919
rect 563842 453859 563902 453919
rect 563962 453859 564022 453919
rect 564082 453859 564142 453919
rect 564202 453859 564262 453919
rect 564322 453859 564382 453919
rect 564442 453859 564502 453919
rect 564562 453859 564622 453919
rect 564682 453859 564742 453919
rect 564802 453859 564862 453919
rect 564922 453859 564982 453919
rect 565042 453859 565102 453919
rect 565162 453859 565222 453919
rect 565282 453859 565342 453919
rect 565402 453859 565462 453919
rect 565522 453859 565582 453919
rect 565642 453859 565702 453919
rect 565762 453859 565822 453919
rect 565882 453859 565942 453919
rect 566002 453859 566062 453919
rect 566122 453859 566182 453919
rect 566242 453859 566302 453919
rect 566362 453859 566422 453919
rect 566482 453859 566542 453919
rect 566602 453859 566662 453919
rect 566722 453859 566782 453919
rect 566842 453859 566902 453919
rect 566962 453859 567022 453919
rect 567082 453859 567142 453919
rect 567202 453859 567262 453919
rect 567322 453859 567382 453919
rect 567442 453859 567502 453919
rect 567562 453859 567622 453919
rect 562102 453799 567622 453859
rect 513703 453756 513937 453773
rect 513703 453556 513720 453756
rect 513920 453556 513937 453756
rect 513703 453539 513937 453556
rect 514137 453756 514371 453773
rect 514137 453556 514154 453756
rect 514354 453556 514371 453756
rect 514137 453539 514371 453556
rect 514571 453756 514805 453773
rect 514571 453556 514588 453756
rect 514788 453556 514805 453756
rect 562102 453739 562222 453799
rect 562282 453739 562342 453799
rect 562402 453739 562462 453799
rect 562522 453739 562582 453799
rect 562642 453739 562702 453799
rect 562762 453739 562822 453799
rect 562882 453739 562942 453799
rect 563002 453739 563062 453799
rect 563122 453739 563182 453799
rect 563242 453739 563302 453799
rect 563362 453739 563422 453799
rect 563482 453739 563542 453799
rect 563602 453739 563662 453799
rect 563722 453739 563782 453799
rect 563842 453739 563902 453799
rect 563962 453739 564022 453799
rect 564082 453739 564142 453799
rect 564202 453739 564262 453799
rect 564322 453739 564382 453799
rect 564442 453739 564502 453799
rect 564562 453739 564622 453799
rect 564682 453739 564742 453799
rect 564802 453739 564862 453799
rect 564922 453739 564982 453799
rect 565042 453739 565102 453799
rect 565162 453739 565222 453799
rect 565282 453739 565342 453799
rect 565402 453739 565462 453799
rect 565522 453739 565582 453799
rect 565642 453739 565702 453799
rect 565762 453739 565822 453799
rect 565882 453739 565942 453799
rect 566002 453739 566062 453799
rect 566122 453739 566182 453799
rect 566242 453739 566302 453799
rect 566362 453739 566422 453799
rect 566482 453739 566542 453799
rect 566602 453739 566662 453799
rect 566722 453739 566782 453799
rect 566842 453739 566902 453799
rect 566962 453739 567022 453799
rect 567082 453739 567142 453799
rect 567202 453739 567262 453799
rect 567322 453739 567382 453799
rect 567442 453739 567502 453799
rect 567562 453739 567622 453799
rect 562102 453679 567622 453739
rect 572272 453934 577792 453994
rect 572272 453874 572332 453934
rect 572392 453874 572452 453934
rect 572512 453874 572572 453934
rect 572632 453874 572692 453934
rect 572752 453874 572812 453934
rect 572872 453874 572932 453934
rect 572992 453874 573052 453934
rect 573112 453874 573172 453934
rect 573232 453874 573292 453934
rect 573352 453874 573412 453934
rect 573472 453874 573532 453934
rect 573592 453874 573652 453934
rect 573712 453874 573772 453934
rect 573832 453874 573892 453934
rect 573952 453874 574012 453934
rect 574072 453874 574132 453934
rect 574192 453874 574252 453934
rect 574312 453874 574372 453934
rect 574432 453874 574492 453934
rect 574552 453874 574612 453934
rect 574672 453874 574732 453934
rect 574792 453874 574852 453934
rect 574912 453874 574972 453934
rect 575032 453874 575092 453934
rect 575152 453874 575212 453934
rect 575272 453874 575332 453934
rect 575392 453874 575452 453934
rect 575512 453874 575572 453934
rect 575632 453874 575692 453934
rect 575752 453874 575812 453934
rect 575872 453874 575932 453934
rect 575992 453874 576052 453934
rect 576112 453874 576172 453934
rect 576232 453874 576292 453934
rect 576352 453874 576412 453934
rect 576472 453874 576532 453934
rect 576592 453874 576652 453934
rect 576712 453874 576772 453934
rect 576832 453874 576892 453934
rect 576952 453874 577012 453934
rect 577072 453874 577132 453934
rect 577192 453874 577252 453934
rect 577312 453874 577372 453934
rect 577432 453874 577492 453934
rect 577552 453874 577612 453934
rect 577672 453874 577792 453934
rect 572272 453814 577792 453874
rect 572272 453754 572332 453814
rect 572392 453754 572452 453814
rect 572512 453754 572572 453814
rect 572632 453754 572692 453814
rect 572752 453754 572812 453814
rect 572872 453754 572932 453814
rect 572992 453754 573052 453814
rect 573112 453754 573172 453814
rect 573232 453754 573292 453814
rect 573352 453754 573412 453814
rect 573472 453754 573532 453814
rect 573592 453754 573652 453814
rect 573712 453754 573772 453814
rect 573832 453754 573892 453814
rect 573952 453754 574012 453814
rect 574072 453754 574132 453814
rect 574192 453754 574252 453814
rect 574312 453754 574372 453814
rect 574432 453754 574492 453814
rect 574552 453754 574612 453814
rect 574672 453754 574732 453814
rect 574792 453754 574852 453814
rect 574912 453754 574972 453814
rect 575032 453754 575092 453814
rect 575152 453754 575212 453814
rect 575272 453754 575332 453814
rect 575392 453754 575452 453814
rect 575512 453754 575572 453814
rect 575632 453754 575692 453814
rect 575752 453754 575812 453814
rect 575872 453754 575932 453814
rect 575992 453754 576052 453814
rect 576112 453754 576172 453814
rect 576232 453754 576292 453814
rect 576352 453754 576412 453814
rect 576472 453754 576532 453814
rect 576592 453754 576652 453814
rect 576712 453754 576772 453814
rect 576832 453754 576892 453814
rect 576952 453754 577012 453814
rect 577072 453754 577132 453814
rect 577192 453754 577252 453814
rect 577312 453754 577372 453814
rect 577432 453754 577492 453814
rect 577552 453754 577612 453814
rect 577672 453754 577792 453814
rect 572272 453694 577792 453754
rect 514571 453539 514805 453556
rect 513703 453322 513937 453339
rect 513703 453122 513720 453322
rect 513920 453122 513937 453322
rect 513703 453105 513937 453122
rect 514137 453322 514371 453339
rect 514137 453122 514154 453322
rect 514354 453122 514371 453322
rect 514137 453105 514371 453122
rect 514571 453322 514805 453339
rect 514571 453122 514588 453322
rect 514788 453122 514805 453322
rect 514571 453105 514805 453122
rect 513703 452888 513937 452905
rect 513703 452688 513720 452888
rect 513920 452688 513937 452888
rect 513703 452671 513937 452688
rect 514137 452888 514371 452905
rect 514137 452688 514154 452888
rect 514354 452688 514371 452888
rect 514137 452671 514371 452688
rect 514571 452888 514805 452905
rect 514571 452688 514588 452888
rect 514788 452688 514805 452888
rect 514571 452671 514805 452688
rect 513703 452454 513937 452471
rect 513703 452254 513720 452454
rect 513920 452254 513937 452454
rect 513703 452237 513937 452254
rect 514137 452454 514371 452471
rect 514137 452254 514154 452454
rect 514354 452254 514371 452454
rect 514137 452237 514371 452254
rect 514571 452454 514805 452471
rect 514571 452254 514588 452454
rect 514788 452254 514805 452454
rect 514571 452237 514805 452254
rect 513703 452020 513937 452037
rect 513703 451820 513720 452020
rect 513920 451820 513937 452020
rect 513703 451803 513937 451820
rect 514137 452020 514371 452037
rect 514137 451820 514154 452020
rect 514354 451820 514371 452020
rect 514137 451803 514371 451820
rect 514571 452020 514805 452037
rect 514571 451820 514588 452020
rect 514788 451820 514805 452020
rect 514571 451803 514805 451820
rect 513703 451586 513937 451603
rect 513703 451386 513720 451586
rect 513920 451386 513937 451586
rect 513703 451369 513937 451386
rect 514137 451586 514371 451603
rect 514137 451386 514154 451586
rect 514354 451386 514371 451586
rect 514137 451369 514371 451386
rect 514571 451586 514805 451603
rect 514571 451386 514588 451586
rect 514788 451386 514805 451586
rect 514571 451369 514805 451386
rect 513703 451152 513937 451169
rect 513703 450952 513720 451152
rect 513920 450952 513937 451152
rect 513703 450935 513937 450952
rect 514137 451152 514371 451169
rect 514137 450952 514154 451152
rect 514354 450952 514371 451152
rect 514137 450935 514371 450952
rect 514571 451152 514805 451169
rect 514571 450952 514588 451152
rect 514788 450952 514805 451152
rect 514571 450935 514805 450952
rect 515390 450880 516622 450886
rect 513703 450718 513937 450735
rect 513703 450518 513720 450718
rect 513920 450518 513937 450718
rect 513703 450501 513937 450518
rect 514137 450718 514371 450735
rect 514137 450518 514154 450718
rect 514354 450518 514371 450718
rect 514137 450501 514371 450518
rect 514571 450718 514805 450735
rect 514571 450518 514588 450718
rect 514788 450518 514805 450718
rect 514571 450501 514805 450518
rect 515390 450322 515396 450880
rect 515954 450322 516196 450880
rect 516616 450322 516622 450880
rect 515396 450316 516622 450322
rect 522126 450880 523358 450886
rect 522126 450322 522132 450880
rect 522690 450322 522932 450880
rect 523352 450322 523358 450880
rect 522126 450316 523358 450322
rect 513703 450284 513937 450301
rect 513703 450084 513720 450284
rect 513920 450084 513937 450284
rect 513703 450067 513937 450084
rect 514137 450284 514371 450301
rect 514137 450084 514154 450284
rect 514354 450084 514371 450284
rect 514137 450067 514371 450084
rect 514571 450284 514805 450301
rect 514571 450084 514588 450284
rect 514788 450084 514805 450284
rect 514571 450067 514805 450084
rect 516190 450062 518222 450068
rect 513703 449850 513937 449867
rect 513703 449650 513720 449850
rect 513920 449650 513937 449850
rect 513703 449633 513937 449650
rect 514137 449850 514371 449867
rect 514137 449650 514154 449850
rect 514354 449650 514371 449850
rect 514137 449633 514371 449650
rect 514571 449850 514805 449867
rect 514571 449650 514588 449850
rect 514788 449650 514805 449850
rect 514571 449633 514805 449650
rect 516190 449504 516196 450062
rect 516616 449504 517658 450062
rect 518216 449504 518222 450062
rect 516190 449498 518222 449504
rect 522926 450062 524158 450068
rect 522926 449504 522932 450062
rect 523352 449504 523594 450062
rect 524152 449504 524158 450062
rect 522926 449498 524158 449504
rect 513703 449416 513937 449433
rect 513703 449216 513720 449416
rect 513920 449216 513937 449416
rect 513703 449199 513937 449216
rect 514137 449416 514371 449433
rect 514137 449216 514154 449416
rect 514354 449216 514371 449416
rect 514137 449199 514371 449216
rect 514571 449416 514805 449433
rect 514571 449216 514588 449416
rect 514788 449216 514805 449416
rect 514571 449199 514805 449216
rect 516190 449244 517422 449250
rect 514571 449016 514805 449033
rect 514571 448816 514588 449016
rect 514788 448816 514805 449016
rect 514571 448799 514805 448816
rect 516190 448686 516196 449244
rect 516616 448686 516858 449244
rect 517416 448686 517422 449244
rect 516190 448680 517422 448686
rect 522926 449244 523358 449250
rect 522926 448686 522932 449244
rect 523352 449238 523358 449244
rect 523352 449232 524958 449238
rect 523352 448686 524394 449232
rect 522926 448680 524394 448686
rect 522944 448674 524394 448680
rect 524952 448674 524958 449232
rect 522944 448668 524958 448674
rect 514571 448616 514805 448633
rect 514571 448416 514588 448616
rect 514788 448416 514805 448616
rect 514571 448399 514805 448416
rect 515390 448426 516622 448432
rect 514571 448216 514805 448233
rect 514571 448016 514588 448216
rect 514788 448016 514805 448216
rect 514571 447999 514805 448016
rect 515390 447868 515396 448426
rect 515954 447868 516196 448426
rect 516616 447868 516622 448426
rect 515396 447862 516622 447868
rect 522126 448426 523358 448432
rect 522126 447868 522132 448426
rect 522690 447868 522932 448426
rect 523352 447868 523358 448426
rect 522126 447862 523358 447868
rect 514571 447816 514805 447833
rect 514571 447616 514588 447816
rect 514788 447616 514805 447816
rect 514571 447599 514805 447616
rect 516190 447608 517422 447614
rect 514571 447416 514805 447433
rect 514571 447216 514588 447416
rect 514788 447216 514805 447416
rect 514571 447199 514805 447216
rect 516190 447050 516196 447608
rect 516616 447050 516858 447608
rect 517416 447050 517422 447608
rect 516190 447044 517422 447050
rect 522926 447608 524958 447614
rect 522926 447050 522932 447608
rect 523352 447050 524394 447608
rect 524952 447050 524958 447608
rect 522926 447044 524958 447050
rect 514571 447016 514805 447033
rect 514571 446816 514588 447016
rect 514788 446816 514805 447016
rect 514571 446799 514805 446816
rect 516190 446790 518222 446796
rect 514571 446616 514805 446633
rect 514571 446416 514588 446616
rect 514788 446416 514805 446616
rect 514571 446399 514805 446416
rect 514571 446216 514805 446233
rect 516190 446232 516196 446790
rect 516616 446232 517658 446790
rect 518216 446232 518222 446790
rect 516190 446226 518222 446232
rect 522926 446790 524158 446796
rect 522926 446232 522932 446790
rect 523352 446232 523594 446790
rect 524152 446232 524158 446790
rect 522926 446226 524158 446232
rect 514571 446016 514588 446216
rect 514788 446016 514805 446216
rect 514571 445999 514805 446016
rect 515390 445972 516622 445978
rect 512112 443648 512134 445636
rect 513286 443648 513294 445636
rect 514571 445816 514805 445833
rect 514571 445616 514588 445816
rect 514788 445616 514805 445816
rect 514571 445599 514805 445616
rect 515390 445414 515396 445972
rect 515954 445414 516196 445972
rect 516616 445414 516622 445972
rect 515396 445408 516622 445414
rect 522126 445972 523358 445978
rect 522126 445414 522132 445972
rect 522690 445414 522932 445972
rect 523352 445414 523358 445972
rect 522126 445408 523358 445414
rect 512112 439882 512228 443648
rect 513212 440324 513294 443648
rect 513542 445232 516584 445238
rect 513542 444540 516066 445232
rect 516584 445154 516622 445160
rect 516616 444596 516622 445154
rect 516584 444590 516622 444596
rect 519926 445154 523358 445160
rect 519926 444596 522932 445154
rect 523352 444596 523358 445154
rect 519926 444590 523358 444596
rect 513542 444536 516584 444540
rect 513542 441666 514072 444536
rect 515318 444534 516584 444536
rect 516190 444336 518222 444342
rect 514571 444216 514805 444233
rect 514571 444016 514588 444216
rect 514788 444016 514805 444216
rect 514571 443999 514805 444016
rect 514571 443816 514805 443833
rect 514571 443616 514588 443816
rect 514788 443616 514805 443816
rect 516190 443778 516196 444336
rect 516616 443778 517658 444336
rect 518216 443778 518222 444336
rect 516190 443772 518222 443778
rect 514571 443599 514805 443616
rect 516190 443518 517422 443524
rect 514571 443416 514805 443433
rect 514571 443216 514588 443416
rect 514788 443216 514805 443416
rect 514571 443199 514805 443216
rect 514571 443016 514805 443033
rect 514571 442816 514588 443016
rect 514788 442816 514805 443016
rect 516190 442960 516196 443518
rect 516616 442960 516858 443518
rect 517416 442960 517422 443518
rect 516190 442954 517422 442960
rect 514571 442799 514805 442816
rect 515390 442700 516622 442706
rect 514571 442616 514805 442633
rect 514571 442416 514588 442616
rect 514788 442416 514805 442616
rect 514571 442399 514805 442416
rect 514571 442216 514805 442233
rect 514571 442016 514588 442216
rect 514788 442016 514805 442216
rect 515390 442142 515396 442700
rect 515954 442142 516196 442700
rect 516616 442142 516622 442700
rect 515390 442136 516622 442142
rect 514571 441999 514805 442016
rect 516190 441882 518222 441888
rect 513542 440732 513548 441666
rect 514066 440732 514072 441666
rect 514571 441816 514805 441833
rect 514571 441616 514588 441816
rect 514788 441616 514805 441816
rect 514571 441599 514805 441616
rect 514571 441416 514805 441433
rect 514571 441216 514588 441416
rect 514788 441216 514805 441416
rect 516190 441324 516196 441882
rect 516616 441324 517658 441882
rect 518216 441324 518222 441882
rect 516190 441318 518222 441324
rect 514571 441199 514805 441216
rect 515918 441142 516622 441148
rect 514571 441016 514805 441033
rect 514571 440816 514588 441016
rect 514788 440816 514805 441016
rect 514571 440799 514805 440816
rect 513542 440726 514072 440732
rect 515918 440450 515924 441142
rect 516616 440450 516622 441142
rect 515918 440444 516622 440450
rect 512112 439632 512836 439882
rect 513286 439632 513294 440324
rect 512112 439612 513294 439632
rect 515924 440324 516622 440330
rect 516616 439632 516622 440324
rect 515924 439626 516622 439632
rect 511228 438814 511534 439504
rect 511822 438814 511828 439504
rect 511228 438808 511828 438814
rect 515918 439506 516622 439512
rect 515918 438814 515924 439506
rect 516616 439446 516622 439506
rect 519926 439446 520496 444590
rect 522926 444336 524158 444342
rect 522926 443778 522932 444336
rect 523352 443778 523594 444336
rect 524152 443778 524158 444336
rect 522926 443772 524158 443778
rect 522926 443518 524958 443524
rect 522926 442960 522932 443518
rect 523352 442960 524394 443518
rect 524952 442960 524958 443518
rect 522926 442954 524958 442960
rect 522126 442700 523358 442706
rect 522126 442142 522132 442700
rect 522690 442142 522932 442700
rect 523352 442142 523358 442700
rect 522126 442136 523358 442142
rect 522926 441882 524158 441888
rect 522926 441324 522932 441882
rect 523352 441324 523594 441882
rect 524152 441324 524158 441882
rect 522926 441318 524158 441324
rect 522926 441064 524388 441070
rect 522926 440506 522932 441064
rect 523352 440506 524394 441064
rect 524952 440506 524958 441064
rect 522926 440500 524958 440506
rect 522126 440246 523358 440252
rect 522126 439688 522132 440246
rect 522690 439688 522932 440246
rect 523352 439688 523358 440246
rect 522126 439682 523358 439688
rect 516616 438876 520496 439446
rect 522926 439428 524158 439434
rect 516616 438814 516622 438876
rect 522926 438870 522932 439428
rect 523352 438870 523594 439428
rect 524152 438870 524158 439428
rect 522926 438864 524158 438870
rect 515918 438808 516622 438814
rect 508800 435508 508868 435560
rect 508920 435508 508972 435560
rect 509024 435508 509076 435560
rect 509128 435508 509180 435560
rect 509232 435508 509284 435560
rect 509336 435508 509388 435560
rect 509440 435508 509504 435560
rect 508800 435456 509504 435508
rect 508800 435404 508868 435456
rect 508920 435404 508972 435456
rect 509024 435404 509076 435456
rect 509128 435404 509180 435456
rect 509232 435404 509284 435456
rect 509336 435404 509388 435456
rect 509440 435404 509504 435456
rect 508800 435352 509504 435404
rect 508800 435300 508868 435352
rect 508920 435300 508972 435352
rect 509024 435300 509076 435352
rect 509128 435300 509180 435352
rect 509232 435300 509284 435352
rect 509336 435300 509388 435352
rect 509440 435300 509504 435352
rect 508800 435248 509504 435300
rect 508800 435196 508868 435248
rect 508920 435196 508972 435248
rect 509024 435196 509076 435248
rect 509128 435196 509180 435248
rect 509232 435196 509284 435248
rect 509336 435196 509388 435248
rect 509440 435196 509504 435248
rect 508800 435144 509504 435196
rect 508800 435092 508868 435144
rect 508920 435092 508972 435144
rect 509024 435092 509076 435144
rect 509128 435092 509180 435144
rect 509232 435092 509284 435144
rect 509336 435092 509388 435144
rect 509440 435092 509504 435144
rect 508800 435040 509504 435092
rect 508800 434988 508868 435040
rect 508920 434988 508972 435040
rect 509024 434988 509076 435040
rect 509128 434988 509180 435040
rect 509232 434988 509284 435040
rect 509336 434988 509388 435040
rect 509440 434988 509504 435040
rect 508800 434936 509504 434988
rect 527604 437540 528664 437580
rect 527604 437440 527638 437540
rect 527738 437440 527862 437540
rect 527962 437440 528086 437540
rect 528186 437440 528310 437540
rect 528410 437440 528534 437540
rect 528634 437440 528664 437540
rect 527604 437316 528664 437440
rect 527604 437216 527638 437316
rect 527738 437216 527862 437316
rect 527962 437216 528086 437316
rect 528186 437216 528310 437316
rect 528410 437216 528534 437316
rect 528634 437216 528664 437316
rect 527604 437092 528664 437216
rect 527604 436992 527638 437092
rect 527738 436992 527862 437092
rect 527962 436992 528086 437092
rect 528186 436992 528310 437092
rect 528410 436992 528534 437092
rect 528634 436992 528664 437092
rect 527604 436868 528664 436992
rect 527604 436768 527638 436868
rect 527738 436768 527862 436868
rect 527962 436768 528086 436868
rect 528186 436768 528310 436868
rect 528410 436768 528534 436868
rect 528634 436768 528664 436868
rect 527604 436644 528664 436768
rect 527604 436544 527638 436644
rect 527738 436544 527862 436644
rect 527962 436544 528086 436644
rect 528186 436544 528310 436644
rect 528410 436544 528534 436644
rect 528634 436544 528664 436644
rect 527604 436420 528664 436544
rect 527604 436320 527638 436420
rect 527738 436320 527862 436420
rect 527962 436320 528086 436420
rect 528186 436320 528310 436420
rect 528410 436320 528534 436420
rect 528634 436320 528664 436420
rect 527604 436196 528664 436320
rect 527604 436096 527638 436196
rect 527738 436096 527862 436196
rect 527962 436096 528086 436196
rect 528186 436096 528310 436196
rect 528410 436096 528534 436196
rect 528634 436096 528664 436196
rect 527604 435972 528664 436096
rect 527604 435872 527638 435972
rect 527738 435872 527862 435972
rect 527962 435872 528086 435972
rect 528186 435872 528310 435972
rect 528410 435872 528534 435972
rect 528634 435872 528664 435972
rect 527604 435748 528664 435872
rect 527604 435648 527638 435748
rect 527738 435648 527862 435748
rect 527962 435648 528086 435748
rect 528186 435648 528310 435748
rect 528410 435648 528534 435748
rect 528634 435648 528664 435748
rect 527604 435524 528664 435648
rect 527604 435424 527638 435524
rect 527738 435424 527862 435524
rect 527962 435424 528086 435524
rect 528186 435424 528310 435524
rect 528410 435424 528534 435524
rect 528634 435424 528664 435524
rect 527604 435300 528664 435424
rect 527604 435200 527638 435300
rect 527738 435200 527862 435300
rect 527962 435200 528086 435300
rect 528186 435200 528310 435300
rect 528410 435200 528534 435300
rect 528634 435200 528664 435300
rect 527604 435076 528664 435200
rect 527604 434976 527638 435076
rect 527738 434976 527862 435076
rect 527962 434976 528086 435076
rect 528186 434976 528310 435076
rect 528410 434976 528534 435076
rect 528634 434976 528664 435076
rect 500384 434752 500418 434852
rect 500518 434752 500642 434852
rect 500742 434752 500866 434852
rect 500966 434752 501090 434852
rect 501190 434752 501314 434852
rect 501414 434752 501444 434852
rect 500384 434628 501444 434752
rect 500384 434528 500418 434628
rect 500518 434528 500642 434628
rect 500742 434528 500866 434628
rect 500966 434528 501090 434628
rect 501190 434528 501314 434628
rect 501414 434528 501444 434628
rect 500384 434404 501444 434528
rect 500384 434304 500418 434404
rect 500518 434304 500642 434404
rect 500742 434304 500866 434404
rect 500966 434304 501090 434404
rect 501190 434304 501314 434404
rect 501414 434304 501444 434404
rect 500384 434180 501444 434304
rect 500384 434080 500418 434180
rect 500518 434080 500642 434180
rect 500742 434080 500866 434180
rect 500966 434080 501090 434180
rect 501190 434080 501314 434180
rect 501414 434080 501444 434180
rect 500384 433956 501444 434080
rect 500384 433856 500418 433956
rect 500518 433856 500642 433956
rect 500742 433856 500866 433956
rect 500966 433856 501090 433956
rect 501190 433856 501314 433956
rect 501414 433856 501444 433956
rect 500384 433732 501444 433856
rect 500384 433632 500418 433732
rect 500518 433632 500642 433732
rect 500742 433632 500866 433732
rect 500966 433632 501090 433732
rect 501190 433632 501314 433732
rect 501414 433632 501444 433732
rect 500384 433508 501444 433632
rect 500384 433408 500418 433508
rect 500518 433408 500642 433508
rect 500742 433408 500866 433508
rect 500966 433408 501090 433508
rect 501190 433408 501314 433508
rect 501414 433408 501444 433508
rect 500384 433284 501444 433408
rect 500384 433184 500418 433284
rect 500518 433184 500642 433284
rect 500742 433184 500866 433284
rect 500966 433184 501090 433284
rect 501190 433184 501314 433284
rect 501414 433184 501444 433284
rect 500384 433060 501444 433184
rect 500384 432960 500418 433060
rect 500518 432960 500642 433060
rect 500742 432960 500866 433060
rect 500966 432960 501090 433060
rect 501190 432960 501314 433060
rect 501414 432960 501444 433060
rect 500384 432836 501444 432960
rect 500384 432736 500418 432836
rect 500518 432736 500642 432836
rect 500742 432736 500866 432836
rect 500966 432736 501090 432836
rect 501190 432736 501314 432836
rect 501414 432736 501444 432836
rect 500384 432612 501444 432736
rect 500384 432512 500418 432612
rect 500518 432512 500642 432612
rect 500742 432512 500866 432612
rect 500966 432512 501090 432612
rect 501190 432512 501314 432612
rect 501414 432512 501444 432612
rect 500384 432388 501444 432512
rect 500384 432288 500418 432388
rect 500518 432288 500642 432388
rect 500742 432288 500866 432388
rect 500966 432288 501090 432388
rect 501190 432288 501314 432388
rect 501414 432288 501444 432388
rect 500384 432164 501444 432288
rect 500384 432064 500418 432164
rect 500518 432064 500642 432164
rect 500742 432064 500866 432164
rect 500966 432064 501090 432164
rect 501190 432064 501314 432164
rect 501414 432064 501444 432164
rect 500384 431940 501444 432064
rect 500384 431840 500418 431940
rect 500518 431840 500642 431940
rect 500742 431840 500866 431940
rect 500966 431840 501090 431940
rect 501190 431840 501314 431940
rect 501414 431840 501444 431940
rect 500384 431716 501444 431840
rect 500384 431616 500418 431716
rect 500518 431616 500642 431716
rect 500742 431616 500866 431716
rect 500966 431616 501090 431716
rect 501190 431616 501314 431716
rect 501414 431616 501444 431716
rect 500384 431492 501444 431616
rect 500384 431392 500418 431492
rect 500518 431392 500642 431492
rect 500742 431392 500866 431492
rect 500966 431392 501090 431492
rect 501190 431392 501314 431492
rect 501414 431392 501444 431492
rect 500384 431268 501444 431392
rect 500384 431168 500418 431268
rect 500518 431168 500642 431268
rect 500742 431168 500866 431268
rect 500966 431168 501090 431268
rect 501190 431168 501314 431268
rect 501414 431168 501444 431268
rect 500384 431044 501444 431168
rect 527604 434852 528664 434976
rect 527604 434752 527638 434852
rect 527738 434752 527862 434852
rect 527962 434752 528086 434852
rect 528186 434752 528310 434852
rect 528410 434752 528534 434852
rect 528634 434752 528664 434852
rect 527604 434628 528664 434752
rect 527604 434528 527638 434628
rect 527738 434528 527862 434628
rect 527962 434528 528086 434628
rect 528186 434528 528310 434628
rect 528410 434528 528534 434628
rect 528634 434528 528664 434628
rect 527604 434404 528664 434528
rect 527604 434304 527638 434404
rect 527738 434304 527862 434404
rect 527962 434304 528086 434404
rect 528186 434304 528310 434404
rect 528410 434304 528534 434404
rect 528634 434304 528664 434404
rect 527604 434180 528664 434304
rect 527604 434080 527638 434180
rect 527738 434080 527862 434180
rect 527962 434080 528086 434180
rect 528186 434080 528310 434180
rect 528410 434080 528534 434180
rect 528634 434080 528664 434180
rect 527604 433956 528664 434080
rect 527604 433856 527638 433956
rect 527738 433856 527862 433956
rect 527962 433856 528086 433956
rect 528186 433856 528310 433956
rect 528410 433856 528534 433956
rect 528634 433856 528664 433956
rect 527604 433732 528664 433856
rect 527604 433632 527638 433732
rect 527738 433632 527862 433732
rect 527962 433632 528086 433732
rect 528186 433632 528310 433732
rect 528410 433632 528534 433732
rect 528634 433632 528664 433732
rect 527604 433508 528664 433632
rect 527604 433408 527638 433508
rect 527738 433408 527862 433508
rect 527962 433408 528086 433508
rect 528186 433408 528310 433508
rect 528410 433408 528534 433508
rect 528634 433408 528664 433508
rect 527604 433284 528664 433408
rect 527604 433184 527638 433284
rect 527738 433184 527862 433284
rect 527962 433184 528086 433284
rect 528186 433184 528310 433284
rect 528410 433184 528534 433284
rect 528634 433184 528664 433284
rect 527604 433060 528664 433184
rect 527604 432960 527638 433060
rect 527738 432960 527862 433060
rect 527962 432960 528086 433060
rect 528186 432960 528310 433060
rect 528410 432960 528534 433060
rect 528634 432960 528664 433060
rect 527604 432836 528664 432960
rect 527604 432736 527638 432836
rect 527738 432736 527862 432836
rect 527962 432736 528086 432836
rect 528186 432736 528310 432836
rect 528410 432736 528534 432836
rect 528634 432736 528664 432836
rect 527604 432612 528664 432736
rect 527604 432512 527638 432612
rect 527738 432512 527862 432612
rect 527962 432512 528086 432612
rect 528186 432512 528310 432612
rect 528410 432512 528534 432612
rect 528634 432512 528664 432612
rect 527604 432388 528664 432512
rect 527604 432288 527638 432388
rect 527738 432288 527862 432388
rect 527962 432288 528086 432388
rect 528186 432288 528310 432388
rect 528410 432288 528534 432388
rect 528634 432288 528664 432388
rect 527604 432164 528664 432288
rect 527604 432064 527638 432164
rect 527738 432064 527862 432164
rect 527962 432064 528086 432164
rect 528186 432064 528310 432164
rect 528410 432064 528534 432164
rect 528634 432064 528664 432164
rect 527604 431940 528664 432064
rect 527604 431840 527638 431940
rect 527738 431840 527862 431940
rect 527962 431840 528086 431940
rect 528186 431840 528310 431940
rect 528410 431840 528534 431940
rect 528634 431840 528664 431940
rect 527604 431716 528664 431840
rect 527604 431616 527638 431716
rect 527738 431616 527862 431716
rect 527962 431616 528086 431716
rect 528186 431616 528310 431716
rect 528410 431616 528534 431716
rect 528634 431616 528664 431716
rect 527604 431492 528664 431616
rect 527604 431392 527638 431492
rect 527738 431392 527862 431492
rect 527962 431392 528086 431492
rect 528186 431392 528310 431492
rect 528410 431392 528534 431492
rect 528634 431392 528664 431492
rect 527604 431268 528664 431392
rect 527604 431168 527638 431268
rect 527738 431168 527862 431268
rect 527962 431168 528086 431268
rect 528186 431168 528310 431268
rect 528410 431168 528534 431268
rect 528634 431168 528664 431268
rect 500384 430944 500418 431044
rect 500518 430944 500642 431044
rect 500742 430944 500866 431044
rect 500966 430944 501090 431044
rect 501190 430944 501314 431044
rect 501414 430944 501444 431044
rect 500384 430920 501444 430944
rect 503900 431026 510526 431056
rect 503900 430926 503920 431026
rect 504020 430926 504144 431026
rect 504244 430926 504368 431026
rect 504468 430926 504592 431026
rect 504692 430926 504816 431026
rect 504916 430926 505040 431026
rect 505140 430926 505264 431026
rect 505364 430926 505488 431026
rect 505588 430926 505712 431026
rect 505812 430926 505936 431026
rect 506036 430926 506160 431026
rect 506260 430926 506384 431026
rect 506484 430926 506608 431026
rect 506708 430926 506832 431026
rect 506932 430926 507056 431026
rect 507156 430926 507280 431026
rect 507380 430926 507504 431026
rect 507604 430926 507728 431026
rect 507828 430926 507952 431026
rect 508052 430926 508176 431026
rect 508276 430926 508400 431026
rect 508500 430926 508624 431026
rect 508724 430926 508848 431026
rect 508948 430926 509072 431026
rect 509172 430926 509296 431026
rect 509396 430926 509520 431026
rect 509620 430926 509744 431026
rect 509844 430926 509968 431026
rect 510068 430926 510192 431026
rect 510292 430926 510416 431026
rect 510516 430926 510526 431026
rect 503900 430802 510526 430926
rect 503900 430702 503920 430802
rect 504020 430702 504144 430802
rect 504244 430702 504368 430802
rect 504468 430702 504592 430802
rect 504692 430702 504816 430802
rect 504916 430702 505040 430802
rect 505140 430702 505264 430802
rect 505364 430702 505488 430802
rect 505588 430702 505712 430802
rect 505812 430702 505936 430802
rect 506036 430702 506160 430802
rect 506260 430702 506384 430802
rect 506484 430702 506608 430802
rect 506708 430702 506832 430802
rect 506932 430702 507056 430802
rect 507156 430702 507280 430802
rect 507380 430702 507504 430802
rect 507604 430702 507728 430802
rect 507828 430702 507952 430802
rect 508052 430702 508176 430802
rect 508276 430702 508400 430802
rect 508500 430702 508624 430802
rect 508724 430702 508848 430802
rect 508948 430702 509072 430802
rect 509172 430702 509296 430802
rect 509396 430702 509520 430802
rect 509620 430702 509744 430802
rect 509844 430702 509968 430802
rect 510068 430702 510192 430802
rect 510292 430702 510416 430802
rect 510516 430702 510526 430802
rect 503900 430578 510526 430702
rect 503900 430478 503920 430578
rect 504020 430478 504144 430578
rect 504244 430478 504368 430578
rect 504468 430478 504592 430578
rect 504692 430478 504816 430578
rect 504916 430478 505040 430578
rect 505140 430478 505264 430578
rect 505364 430478 505488 430578
rect 505588 430478 505712 430578
rect 505812 430478 505936 430578
rect 506036 430478 506160 430578
rect 506260 430478 506384 430578
rect 506484 430478 506608 430578
rect 506708 430478 506832 430578
rect 506932 430478 507056 430578
rect 507156 430478 507280 430578
rect 507380 430478 507504 430578
rect 507604 430478 507728 430578
rect 507828 430478 507952 430578
rect 508052 430478 508176 430578
rect 508276 430478 508400 430578
rect 508500 430478 508624 430578
rect 508724 430478 508848 430578
rect 508948 430478 509072 430578
rect 509172 430478 509296 430578
rect 509396 430478 509520 430578
rect 509620 430478 509744 430578
rect 509844 430478 509968 430578
rect 510068 430478 510192 430578
rect 510292 430478 510416 430578
rect 510516 430478 510526 430578
rect 503900 430354 510526 430478
rect 503900 430254 503920 430354
rect 504020 430254 504144 430354
rect 504244 430254 504368 430354
rect 504468 430254 504592 430354
rect 504692 430254 504816 430354
rect 504916 430254 505040 430354
rect 505140 430254 505264 430354
rect 505364 430254 505488 430354
rect 505588 430254 505712 430354
rect 505812 430254 505936 430354
rect 506036 430254 506160 430354
rect 506260 430254 506384 430354
rect 506484 430254 506608 430354
rect 506708 430254 506832 430354
rect 506932 430254 507056 430354
rect 507156 430254 507280 430354
rect 507380 430254 507504 430354
rect 507604 430254 507728 430354
rect 507828 430254 507952 430354
rect 508052 430254 508176 430354
rect 508276 430254 508400 430354
rect 508500 430254 508624 430354
rect 508724 430254 508848 430354
rect 508948 430254 509072 430354
rect 509172 430254 509296 430354
rect 509396 430254 509520 430354
rect 509620 430254 509744 430354
rect 509844 430254 509968 430354
rect 510068 430254 510192 430354
rect 510292 430254 510416 430354
rect 510516 430254 510526 430354
rect 503900 430130 510526 430254
rect 503900 430030 503920 430130
rect 504020 430030 504144 430130
rect 504244 430030 504368 430130
rect 504468 430030 504592 430130
rect 504692 430030 504816 430130
rect 504916 430030 505040 430130
rect 505140 430030 505264 430130
rect 505364 430030 505488 430130
rect 505588 430030 505712 430130
rect 505812 430030 505936 430130
rect 506036 430030 506160 430130
rect 506260 430030 506384 430130
rect 506484 430030 506608 430130
rect 506708 430030 506832 430130
rect 506932 430030 507056 430130
rect 507156 430030 507280 430130
rect 507380 430030 507504 430130
rect 507604 430030 507728 430130
rect 507828 430030 507952 430130
rect 508052 430030 508176 430130
rect 508276 430030 508400 430130
rect 508500 430030 508624 430130
rect 508724 430030 508848 430130
rect 508948 430030 509072 430130
rect 509172 430030 509296 430130
rect 509396 430030 509520 430130
rect 509620 430030 509744 430130
rect 509844 430030 509968 430130
rect 510068 430030 510192 430130
rect 510292 430030 510416 430130
rect 510516 430030 510526 430130
rect 503900 429998 510526 430030
rect 517280 431026 523940 431056
rect 517280 430926 517320 431026
rect 517420 430926 517544 431026
rect 517644 430926 517768 431026
rect 517868 430926 517992 431026
rect 518092 430926 518216 431026
rect 518316 430926 518440 431026
rect 518540 430926 518664 431026
rect 518764 430926 518888 431026
rect 518988 430926 519112 431026
rect 519212 430926 519336 431026
rect 519436 430926 519560 431026
rect 519660 430926 519784 431026
rect 519884 430926 520008 431026
rect 520108 430926 520232 431026
rect 520332 430926 520456 431026
rect 520556 430926 520680 431026
rect 520780 430926 520904 431026
rect 521004 430926 521128 431026
rect 521228 430926 521352 431026
rect 521452 430926 521576 431026
rect 521676 430926 521800 431026
rect 521900 430926 522024 431026
rect 522124 430926 522248 431026
rect 522348 430926 522472 431026
rect 522572 430926 522696 431026
rect 522796 430926 522920 431026
rect 523020 430926 523144 431026
rect 523244 430926 523368 431026
rect 523468 430926 523592 431026
rect 523692 430926 523816 431026
rect 523916 430926 523940 431026
rect 517280 430802 523940 430926
rect 527604 431044 528664 431168
rect 527604 430944 527638 431044
rect 527738 430944 527862 431044
rect 527962 430944 528086 431044
rect 528186 430944 528310 431044
rect 528410 430944 528534 431044
rect 528634 430944 528664 431044
rect 527604 430920 528664 430944
rect 517280 430702 517320 430802
rect 517420 430702 517544 430802
rect 517644 430702 517768 430802
rect 517868 430702 517992 430802
rect 518092 430702 518216 430802
rect 518316 430702 518440 430802
rect 518540 430702 518664 430802
rect 518764 430702 518888 430802
rect 518988 430702 519112 430802
rect 519212 430702 519336 430802
rect 519436 430702 519560 430802
rect 519660 430702 519784 430802
rect 519884 430702 520008 430802
rect 520108 430702 520232 430802
rect 520332 430702 520456 430802
rect 520556 430702 520680 430802
rect 520780 430702 520904 430802
rect 521004 430702 521128 430802
rect 521228 430702 521352 430802
rect 521452 430702 521576 430802
rect 521676 430702 521800 430802
rect 521900 430702 522024 430802
rect 522124 430702 522248 430802
rect 522348 430702 522472 430802
rect 522572 430702 522696 430802
rect 522796 430702 522920 430802
rect 523020 430702 523144 430802
rect 523244 430702 523368 430802
rect 523468 430702 523592 430802
rect 523692 430702 523816 430802
rect 523916 430702 523940 430802
rect 517280 430578 523940 430702
rect 517280 430478 517320 430578
rect 517420 430478 517544 430578
rect 517644 430478 517768 430578
rect 517868 430478 517992 430578
rect 518092 430478 518216 430578
rect 518316 430478 518440 430578
rect 518540 430478 518664 430578
rect 518764 430478 518888 430578
rect 518988 430478 519112 430578
rect 519212 430478 519336 430578
rect 519436 430478 519560 430578
rect 519660 430478 519784 430578
rect 519884 430478 520008 430578
rect 520108 430478 520232 430578
rect 520332 430478 520456 430578
rect 520556 430478 520680 430578
rect 520780 430478 520904 430578
rect 521004 430478 521128 430578
rect 521228 430478 521352 430578
rect 521452 430478 521576 430578
rect 521676 430478 521800 430578
rect 521900 430478 522024 430578
rect 522124 430478 522248 430578
rect 522348 430478 522472 430578
rect 522572 430478 522696 430578
rect 522796 430478 522920 430578
rect 523020 430478 523144 430578
rect 523244 430478 523368 430578
rect 523468 430478 523592 430578
rect 523692 430478 523816 430578
rect 523916 430478 523940 430578
rect 517280 430354 523940 430478
rect 517280 430254 517320 430354
rect 517420 430254 517544 430354
rect 517644 430254 517768 430354
rect 517868 430254 517992 430354
rect 518092 430254 518216 430354
rect 518316 430254 518440 430354
rect 518540 430254 518664 430354
rect 518764 430254 518888 430354
rect 518988 430254 519112 430354
rect 519212 430254 519336 430354
rect 519436 430254 519560 430354
rect 519660 430254 519784 430354
rect 519884 430254 520008 430354
rect 520108 430254 520232 430354
rect 520332 430254 520456 430354
rect 520556 430254 520680 430354
rect 520780 430254 520904 430354
rect 521004 430254 521128 430354
rect 521228 430254 521352 430354
rect 521452 430254 521576 430354
rect 521676 430254 521800 430354
rect 521900 430254 522024 430354
rect 522124 430254 522248 430354
rect 522348 430254 522472 430354
rect 522572 430254 522696 430354
rect 522796 430254 522920 430354
rect 523020 430254 523144 430354
rect 523244 430254 523368 430354
rect 523468 430254 523592 430354
rect 523692 430254 523816 430354
rect 523916 430254 523940 430354
rect 517280 430130 523940 430254
rect 517280 430030 517320 430130
rect 517420 430030 517544 430130
rect 517644 430030 517768 430130
rect 517868 430030 517992 430130
rect 518092 430030 518216 430130
rect 518316 430030 518440 430130
rect 518540 430030 518664 430130
rect 518764 430030 518888 430130
rect 518988 430030 519112 430130
rect 519212 430030 519336 430130
rect 519436 430030 519560 430130
rect 519660 430030 519784 430130
rect 519884 430030 520008 430130
rect 520108 430030 520232 430130
rect 520332 430030 520456 430130
rect 520556 430030 520680 430130
rect 520780 430030 520904 430130
rect 521004 430030 521128 430130
rect 521228 430030 521352 430130
rect 521452 430030 521576 430130
rect 521676 430030 521800 430130
rect 521900 430030 522024 430130
rect 522124 430030 522248 430130
rect 522348 430030 522472 430130
rect 522572 430030 522696 430130
rect 522796 430030 522920 430130
rect 523020 430030 523144 430130
rect 523244 430030 523368 430130
rect 523468 430030 523592 430130
rect 523692 430030 523816 430130
rect 523916 430030 523940 430130
rect 517280 429996 523940 430030
rect 524 -800 636 480
rect 1706 -800 1818 480
rect 2888 -800 3000 480
rect 4070 -800 4182 480
rect 5252 -800 5364 480
rect 6434 -800 6546 480
rect 7616 -800 7728 480
rect 8798 -800 8910 480
rect 9980 -800 10092 480
rect 11162 -800 11274 480
rect 12344 -800 12456 480
rect 13526 -800 13638 480
rect 14708 -800 14820 480
rect 15890 -800 16002 480
rect 17072 -800 17184 480
rect 18254 -800 18366 480
rect 19436 -800 19548 480
rect 20618 -800 20730 480
rect 21800 -800 21912 480
rect 22982 -800 23094 480
rect 24164 -800 24276 480
rect 25346 -800 25458 480
rect 26528 -800 26640 480
rect 27710 -800 27822 480
rect 28892 -800 29004 480
rect 30074 -800 30186 480
rect 31256 -800 31368 480
rect 32438 -800 32550 480
rect 33620 -800 33732 480
rect 34802 -800 34914 480
rect 35984 -800 36096 480
rect 37166 -800 37278 480
rect 38348 -800 38460 480
rect 39530 -800 39642 480
rect 40712 -800 40824 480
rect 41894 -800 42006 480
rect 43076 -800 43188 480
rect 44258 -800 44370 480
rect 45440 -800 45552 480
rect 46622 -800 46734 480
rect 47804 -800 47916 480
rect 48986 -800 49098 480
rect 50168 -800 50280 480
rect 51350 -800 51462 480
rect 52532 -800 52644 480
rect 53714 -800 53826 480
rect 54896 -800 55008 480
rect 56078 -800 56190 480
rect 57260 -800 57372 480
rect 58442 -800 58554 480
rect 59624 -800 59736 480
rect 60806 -800 60918 480
rect 61988 -800 62100 480
rect 63170 -800 63282 480
rect 64352 -800 64464 480
rect 65534 -800 65646 480
rect 66716 -800 66828 480
rect 67898 -800 68010 480
rect 69080 -800 69192 480
rect 70262 -800 70374 480
rect 71444 -800 71556 480
rect 72626 -800 72738 480
rect 73808 -800 73920 480
rect 74990 -800 75102 480
rect 76172 -800 76284 480
rect 77354 -800 77466 480
rect 78536 -800 78648 480
rect 79718 -800 79830 480
rect 80900 -800 81012 480
rect 82082 -800 82194 480
rect 83264 -800 83376 480
rect 84446 -800 84558 480
rect 85628 -800 85740 480
rect 86810 -800 86922 480
rect 87992 -800 88104 480
rect 89174 -800 89286 480
rect 90356 -800 90468 480
rect 91538 -800 91650 480
rect 92720 -800 92832 480
rect 93902 -800 94014 480
rect 95084 -800 95196 480
rect 96266 -800 96378 480
rect 97448 -800 97560 480
rect 98630 -800 98742 480
rect 99812 -800 99924 480
rect 100994 -800 101106 480
rect 102176 -800 102288 480
rect 103358 -800 103470 480
rect 104540 -800 104652 480
rect 105722 -800 105834 480
rect 106904 -800 107016 480
rect 108086 -800 108198 480
rect 109268 -800 109380 480
rect 110450 -800 110562 480
rect 111632 -800 111744 480
rect 112814 -800 112926 480
rect 113996 -800 114108 480
rect 115178 -800 115290 480
rect 116360 -800 116472 480
rect 117542 -800 117654 480
rect 118724 -800 118836 480
rect 119906 -800 120018 480
rect 121088 -800 121200 480
rect 122270 -800 122382 480
rect 123452 -800 123564 480
rect 124634 -800 124746 480
rect 125816 -800 125928 480
rect 126998 -800 127110 480
rect 128180 -800 128292 480
rect 129362 -800 129474 480
rect 130544 -800 130656 480
rect 131726 -800 131838 480
rect 132908 -800 133020 480
rect 134090 -800 134202 480
rect 135272 -800 135384 480
rect 136454 -800 136566 480
rect 137636 -800 137748 480
rect 138818 -800 138930 480
rect 140000 -800 140112 480
rect 141182 -800 141294 480
rect 142364 -800 142476 480
rect 143546 -800 143658 480
rect 144728 -800 144840 480
rect 145910 -800 146022 480
rect 147092 -800 147204 480
rect 148274 -800 148386 480
rect 149456 -800 149568 480
rect 150638 -800 150750 480
rect 151820 -800 151932 480
rect 153002 -800 153114 480
rect 154184 -800 154296 480
rect 155366 -800 155478 480
rect 156548 -800 156660 480
rect 157730 -800 157842 480
rect 158912 -800 159024 480
rect 160094 -800 160206 480
rect 161276 -800 161388 480
rect 162458 -800 162570 480
rect 163640 -800 163752 480
rect 164822 -800 164934 480
rect 166004 -800 166116 480
rect 167186 -800 167298 480
rect 168368 -800 168480 480
rect 169550 -800 169662 480
rect 170732 -800 170844 480
rect 171914 -800 172026 480
rect 173096 -800 173208 480
rect 174278 -800 174390 480
rect 175460 -800 175572 480
rect 176642 -800 176754 480
rect 177824 -800 177936 480
rect 179006 -800 179118 480
rect 180188 -800 180300 480
rect 181370 -800 181482 480
rect 182552 -800 182664 480
rect 183734 -800 183846 480
rect 184916 -800 185028 480
rect 186098 -800 186210 480
rect 187280 -800 187392 480
rect 188462 -800 188574 480
rect 189644 -800 189756 480
rect 190826 -800 190938 480
rect 192008 -800 192120 480
rect 193190 -800 193302 480
rect 194372 -800 194484 480
rect 195554 -800 195666 480
rect 196736 -800 196848 480
rect 197918 -800 198030 480
rect 199100 -800 199212 480
rect 200282 -800 200394 480
rect 201464 -800 201576 480
rect 202646 -800 202758 480
rect 203828 -800 203940 480
rect 205010 -800 205122 480
rect 206192 -800 206304 480
rect 207374 -800 207486 480
rect 208556 -800 208668 480
rect 209738 -800 209850 480
rect 210920 -800 211032 480
rect 212102 -800 212214 480
rect 213284 -800 213396 480
rect 214466 -800 214578 480
rect 215648 -800 215760 480
rect 216830 -800 216942 480
rect 218012 -800 218124 480
rect 219194 -800 219306 480
rect 220376 -800 220488 480
rect 221558 -800 221670 480
rect 222740 -800 222852 480
rect 223922 -800 224034 480
rect 225104 -800 225216 480
rect 226286 -800 226398 480
rect 227468 -800 227580 480
rect 228650 -800 228762 480
rect 229832 -800 229944 480
rect 231014 -800 231126 480
rect 232196 -800 232308 480
rect 233378 -800 233490 480
rect 234560 -800 234672 480
rect 235742 -800 235854 480
rect 236924 -800 237036 480
rect 238106 -800 238218 480
rect 239288 -800 239400 480
rect 240470 -800 240582 480
rect 241652 -800 241764 480
rect 242834 -800 242946 480
rect 244016 -800 244128 480
rect 245198 -800 245310 480
rect 246380 -800 246492 480
rect 247562 -800 247674 480
rect 248744 -800 248856 480
rect 249926 -800 250038 480
rect 251108 -800 251220 480
rect 252290 -800 252402 480
rect 253472 -800 253584 480
rect 254654 -800 254766 480
rect 255836 -800 255948 480
rect 257018 -800 257130 480
rect 258200 -800 258312 480
rect 259382 -800 259494 480
rect 260564 -800 260676 480
rect 261746 -800 261858 480
rect 262928 -800 263040 480
rect 264110 -800 264222 480
rect 265292 -800 265404 480
rect 266474 -800 266586 480
rect 267656 -800 267768 480
rect 268838 -800 268950 480
rect 270020 -800 270132 480
rect 271202 -800 271314 480
rect 272384 -800 272496 480
rect 273566 -800 273678 480
rect 274748 -800 274860 480
rect 275930 -800 276042 480
rect 277112 -800 277224 480
rect 278294 -800 278406 480
rect 279476 -800 279588 480
rect 280658 -800 280770 480
rect 281840 -800 281952 480
rect 283022 -800 283134 480
rect 284204 -800 284316 480
rect 285386 -800 285498 480
rect 286568 -800 286680 480
rect 287750 -800 287862 480
rect 288932 -800 289044 480
rect 290114 -800 290226 480
rect 291296 -800 291408 480
rect 292478 -800 292590 480
rect 293660 -800 293772 480
rect 294842 -800 294954 480
rect 296024 -800 296136 480
rect 297206 -800 297318 480
rect 298388 -800 298500 480
rect 299570 -800 299682 480
rect 300752 -800 300864 480
rect 301934 -800 302046 480
rect 303116 -800 303228 480
rect 304298 -800 304410 480
rect 305480 -800 305592 480
rect 306662 -800 306774 480
rect 307844 -800 307956 480
rect 309026 -800 309138 480
rect 310208 -800 310320 480
rect 311390 -800 311502 480
rect 312572 -800 312684 480
rect 313754 -800 313866 480
rect 314936 -800 315048 480
rect 316118 -800 316230 480
rect 317300 -800 317412 480
rect 318482 -800 318594 480
rect 319664 -800 319776 480
rect 320846 -800 320958 480
rect 322028 -800 322140 480
rect 323210 -800 323322 480
rect 324392 -800 324504 480
rect 325574 -800 325686 480
rect 326756 -800 326868 480
rect 327938 -800 328050 480
rect 329120 -800 329232 480
rect 330302 -800 330414 480
rect 331484 -800 331596 480
rect 332666 -800 332778 480
rect 333848 -800 333960 480
rect 335030 -800 335142 480
rect 336212 -800 336324 480
rect 337394 -800 337506 480
rect 338576 -800 338688 480
rect 339758 -800 339870 480
rect 340940 -800 341052 480
rect 342122 -800 342234 480
rect 343304 -800 343416 480
rect 344486 -800 344598 480
rect 345668 -800 345780 480
rect 346850 -800 346962 480
rect 348032 -800 348144 480
rect 349214 -800 349326 480
rect 350396 -800 350508 480
rect 351578 -800 351690 480
rect 352760 -800 352872 480
rect 353942 -800 354054 480
rect 355124 -800 355236 480
rect 356306 -800 356418 480
rect 357488 -800 357600 480
rect 358670 -800 358782 480
rect 359852 -800 359964 480
rect 361034 -800 361146 480
rect 362216 -800 362328 480
rect 363398 -800 363510 480
rect 364580 -800 364692 480
rect 365762 -800 365874 480
rect 366944 -800 367056 480
rect 368126 -800 368238 480
rect 369308 -800 369420 480
rect 370490 -800 370602 480
rect 371672 -800 371784 480
rect 372854 -800 372966 480
rect 374036 -800 374148 480
rect 375218 -800 375330 480
rect 376400 -800 376512 480
rect 377582 -800 377694 480
rect 378764 -800 378876 480
rect 379946 -800 380058 480
rect 381128 -800 381240 480
rect 382310 -800 382422 480
rect 383492 -800 383604 480
rect 384674 -800 384786 480
rect 385856 -800 385968 480
rect 387038 -800 387150 480
rect 388220 -800 388332 480
rect 389402 -800 389514 480
rect 390584 -800 390696 480
rect 391766 -800 391878 480
rect 392948 -800 393060 480
rect 394130 -800 394242 480
rect 395312 -800 395424 480
rect 396494 -800 396606 480
rect 397676 -800 397788 480
rect 398858 -800 398970 480
rect 400040 -800 400152 480
rect 401222 -800 401334 480
rect 402404 -800 402516 480
rect 403586 -800 403698 480
rect 404768 -800 404880 480
rect 405950 -800 406062 480
rect 407132 -800 407244 480
rect 408314 -800 408426 480
rect 409496 -800 409608 480
rect 410678 -800 410790 480
rect 411860 -800 411972 480
rect 413042 -800 413154 480
rect 414224 -800 414336 480
rect 415406 -800 415518 480
rect 416588 -800 416700 480
rect 417770 -800 417882 480
rect 418952 -800 419064 480
rect 420134 -800 420246 480
rect 421316 -800 421428 480
rect 422498 -800 422610 480
rect 423680 -800 423792 480
rect 424862 -800 424974 480
rect 426044 -800 426156 480
rect 427226 -800 427338 480
rect 428408 -800 428520 480
rect 429590 -800 429702 480
rect 430772 -800 430884 480
rect 431954 -800 432066 480
rect 433136 -800 433248 480
rect 434318 -800 434430 480
rect 435500 -800 435612 480
rect 436682 -800 436794 480
rect 437864 -800 437976 480
rect 439046 -800 439158 480
rect 440228 -800 440340 480
rect 441410 -800 441522 480
rect 442592 -800 442704 480
rect 443774 -800 443886 480
rect 444956 -800 445068 480
rect 446138 -800 446250 480
rect 447320 -800 447432 480
rect 448502 -800 448614 480
rect 449684 -800 449796 480
rect 450866 -800 450978 480
rect 452048 -800 452160 480
rect 453230 -800 453342 480
rect 454412 -800 454524 480
rect 455594 -800 455706 480
rect 456776 -800 456888 480
rect 457958 -800 458070 480
rect 459140 -800 459252 480
rect 460322 -800 460434 480
rect 461504 -800 461616 480
rect 462686 -800 462798 480
rect 463868 -800 463980 480
rect 465050 -800 465162 480
rect 466232 -800 466344 480
rect 467414 -800 467526 480
rect 468596 -800 468708 480
rect 469778 -800 469890 480
rect 470960 -800 471072 480
rect 472142 -800 472254 480
rect 473324 -800 473436 480
rect 474506 -800 474618 480
rect 475688 -800 475800 480
rect 476870 -800 476982 480
rect 478052 -800 478164 480
rect 479234 -800 479346 480
rect 480416 -800 480528 480
rect 481598 -800 481710 480
rect 482780 -800 482892 480
rect 483962 -800 484074 480
rect 485144 -800 485256 480
rect 486326 -800 486438 480
rect 487508 -800 487620 480
rect 488690 -800 488802 480
rect 489872 -800 489984 480
rect 491054 -800 491166 480
rect 492236 -800 492348 480
rect 493418 -800 493530 480
rect 494600 -800 494712 480
rect 495782 -800 495894 480
rect 496964 -800 497076 480
rect 498146 -800 498258 480
rect 499328 -800 499440 480
rect 500510 -800 500622 480
rect 501692 -800 501804 480
rect 502874 -800 502986 480
rect 504056 -800 504168 480
rect 505238 -800 505350 480
rect 506420 -800 506532 480
rect 507602 -800 507714 480
rect 508784 -800 508896 480
rect 509966 -800 510078 480
rect 511148 -800 511260 480
rect 512330 -800 512442 480
rect 513512 -800 513624 480
rect 514694 -800 514806 480
rect 515876 -800 515988 480
rect 517058 -800 517170 480
rect 518240 -800 518352 480
rect 519422 -800 519534 480
rect 520604 -800 520716 480
rect 521786 -800 521898 480
rect 522968 -800 523080 480
rect 524150 -800 524262 480
rect 525332 -800 525444 480
rect 526514 -800 526626 480
rect 527696 -800 527808 480
rect 528878 -800 528990 480
rect 530060 -800 530172 480
rect 531242 -800 531354 480
rect 532424 -800 532536 480
rect 533606 -800 533718 480
rect 534788 -800 534900 480
rect 535970 -800 536082 480
rect 537152 -800 537264 480
rect 538334 -800 538446 480
rect 539516 -800 539628 480
rect 540698 -800 540810 480
rect 541880 -800 541992 480
rect 543062 -800 543174 480
rect 544244 -800 544356 480
rect 545426 -800 545538 480
rect 546608 -800 546720 480
rect 547790 -800 547902 480
rect 548972 -800 549084 480
rect 550154 -800 550266 480
rect 551336 -800 551448 480
rect 552518 -800 552630 480
rect 553700 -800 553812 480
rect 554882 -800 554994 480
rect 556064 -800 556176 480
rect 557246 -800 557358 480
rect 558428 -800 558540 480
rect 559610 -800 559722 480
rect 560792 -800 560904 480
rect 561974 -800 562086 480
rect 563156 -800 563268 480
rect 564338 -800 564450 480
rect 565520 -800 565632 480
rect 566702 -800 566814 480
rect 567884 -800 567996 480
rect 569066 -800 569178 480
rect 570248 -800 570360 480
rect 571430 -800 571542 480
rect 572612 -800 572724 480
rect 573794 -800 573906 480
rect 574976 -800 575088 480
rect 576158 -800 576270 480
rect 577340 -800 577452 480
rect 578522 -800 578634 480
rect 579704 -800 579816 480
rect 580886 -800 580998 480
rect 582068 -800 582180 480
rect 583250 -800 583362 480
<< via2 >>
rect 562480 495662 562560 495742
rect 562640 495662 562720 495742
rect 562800 495662 562880 495742
rect 562960 495662 563040 495742
rect 563120 495662 563200 495742
rect 563280 495662 563360 495742
rect 563440 495662 563520 495742
rect 563600 495662 563680 495742
rect 563760 495662 563840 495742
rect 563920 495662 564000 495742
rect 564080 495662 564160 495742
rect 564240 495662 564320 495742
rect 564400 495662 564480 495742
rect 564560 495662 564640 495742
rect 564720 495662 564800 495742
rect 564880 495662 564960 495742
rect 565040 495662 565120 495742
rect 565200 495662 565280 495742
rect 565360 495662 565440 495742
rect 565520 495662 565600 495742
rect 565680 495662 565760 495742
rect 565840 495662 565920 495742
rect 566000 495662 566080 495742
rect 566160 495662 566240 495742
rect 566320 495662 566400 495742
rect 566480 495662 566560 495742
rect 566640 495662 566720 495742
rect 566800 495662 566880 495742
rect 566960 495662 567040 495742
rect 567120 495662 567200 495742
rect 567280 495662 567360 495742
rect 562480 495502 562560 495582
rect 562640 495502 562720 495582
rect 562800 495502 562880 495582
rect 562960 495502 563040 495582
rect 563120 495502 563200 495582
rect 563280 495502 563360 495582
rect 563440 495502 563520 495582
rect 563600 495502 563680 495582
rect 563760 495502 563840 495582
rect 563920 495502 564000 495582
rect 564080 495502 564160 495582
rect 564240 495502 564320 495582
rect 564400 495502 564480 495582
rect 564560 495502 564640 495582
rect 564720 495502 564800 495582
rect 564880 495502 564960 495582
rect 565040 495502 565120 495582
rect 565200 495502 565280 495582
rect 565360 495502 565440 495582
rect 565520 495502 565600 495582
rect 565680 495502 565760 495582
rect 565840 495502 565920 495582
rect 566000 495502 566080 495582
rect 566160 495502 566240 495582
rect 566320 495502 566400 495582
rect 566480 495502 566560 495582
rect 566640 495502 566720 495582
rect 566800 495502 566880 495582
rect 566960 495502 567040 495582
rect 567120 495502 567200 495582
rect 567280 495502 567360 495582
rect 572640 495662 572720 495742
rect 572800 495662 572880 495742
rect 572960 495662 573040 495742
rect 573120 495662 573200 495742
rect 573280 495662 573360 495742
rect 573440 495662 573520 495742
rect 573600 495662 573680 495742
rect 573760 495662 573840 495742
rect 573920 495662 574000 495742
rect 574080 495662 574160 495742
rect 574240 495662 574320 495742
rect 574400 495662 574480 495742
rect 574560 495662 574640 495742
rect 574720 495662 574800 495742
rect 574880 495662 574960 495742
rect 575040 495662 575120 495742
rect 575200 495662 575280 495742
rect 575360 495662 575440 495742
rect 575520 495662 575600 495742
rect 575680 495662 575760 495742
rect 575840 495662 575920 495742
rect 576000 495662 576080 495742
rect 576160 495662 576240 495742
rect 576320 495662 576400 495742
rect 576480 495662 576560 495742
rect 576640 495662 576720 495742
rect 576800 495662 576880 495742
rect 576960 495662 577040 495742
rect 577120 495662 577200 495742
rect 577280 495662 577360 495742
rect 577440 495662 577520 495742
rect 572640 495502 572720 495582
rect 572800 495502 572880 495582
rect 572960 495502 573040 495582
rect 573120 495502 573200 495582
rect 573280 495502 573360 495582
rect 573440 495502 573520 495582
rect 573600 495502 573680 495582
rect 573760 495502 573840 495582
rect 573920 495502 574000 495582
rect 574080 495502 574160 495582
rect 574240 495502 574320 495582
rect 574400 495502 574480 495582
rect 574560 495502 574640 495582
rect 574720 495502 574800 495582
rect 574880 495502 574960 495582
rect 575040 495502 575120 495582
rect 575200 495502 575280 495582
rect 575360 495502 575440 495582
rect 575520 495502 575600 495582
rect 575680 495502 575760 495582
rect 575840 495502 575920 495582
rect 576000 495502 576080 495582
rect 576160 495502 576240 495582
rect 576320 495502 576400 495582
rect 576480 495502 576560 495582
rect 576640 495502 576720 495582
rect 576800 495502 576880 495582
rect 576960 495502 577040 495582
rect 577120 495502 577200 495582
rect 577280 495502 577360 495582
rect 577440 495502 577520 495582
rect 562222 494161 562282 494221
rect 562342 494161 562402 494221
rect 562462 494161 562522 494221
rect 562582 494161 562642 494221
rect 562702 494161 562762 494221
rect 562822 494161 562882 494221
rect 562942 494161 563002 494221
rect 563062 494161 563122 494221
rect 563182 494161 563242 494221
rect 563302 494161 563362 494221
rect 563422 494161 563482 494221
rect 563542 494161 563602 494221
rect 563662 494161 563722 494221
rect 563782 494161 563842 494221
rect 563902 494161 563962 494221
rect 564022 494161 564082 494221
rect 564142 494161 564202 494221
rect 564262 494161 564322 494221
rect 564382 494161 564442 494221
rect 564502 494161 564562 494221
rect 564622 494161 564682 494221
rect 564742 494161 564802 494221
rect 564862 494161 564922 494221
rect 564982 494161 565042 494221
rect 565102 494161 565162 494221
rect 565222 494161 565282 494221
rect 565342 494161 565402 494221
rect 565462 494161 565522 494221
rect 565582 494161 565642 494221
rect 565702 494161 565762 494221
rect 565822 494161 565882 494221
rect 565942 494161 566002 494221
rect 566062 494161 566122 494221
rect 566182 494161 566242 494221
rect 566302 494161 566362 494221
rect 566422 494161 566482 494221
rect 566542 494161 566602 494221
rect 566662 494161 566722 494221
rect 566782 494161 566842 494221
rect 566902 494161 566962 494221
rect 567022 494161 567082 494221
rect 567142 494161 567202 494221
rect 567262 494161 567322 494221
rect 567382 494161 567442 494221
rect 567502 494161 567562 494221
rect 562222 494041 562282 494101
rect 562342 494041 562402 494101
rect 562462 494041 562522 494101
rect 562582 494041 562642 494101
rect 562702 494041 562762 494101
rect 562822 494041 562882 494101
rect 562942 494041 563002 494101
rect 563062 494041 563122 494101
rect 563182 494041 563242 494101
rect 563302 494041 563362 494101
rect 563422 494041 563482 494101
rect 563542 494041 563602 494101
rect 563662 494041 563722 494101
rect 563782 494041 563842 494101
rect 563902 494041 563962 494101
rect 564022 494041 564082 494101
rect 564142 494041 564202 494101
rect 564262 494041 564322 494101
rect 564382 494041 564442 494101
rect 564502 494041 564562 494101
rect 564622 494041 564682 494101
rect 564742 494041 564802 494101
rect 564862 494041 564922 494101
rect 564982 494041 565042 494101
rect 565102 494041 565162 494101
rect 565222 494041 565282 494101
rect 565342 494041 565402 494101
rect 565462 494041 565522 494101
rect 565582 494041 565642 494101
rect 565702 494041 565762 494101
rect 565822 494041 565882 494101
rect 565942 494041 566002 494101
rect 566062 494041 566122 494101
rect 566182 494041 566242 494101
rect 566302 494041 566362 494101
rect 566422 494041 566482 494101
rect 566542 494041 566602 494101
rect 566662 494041 566722 494101
rect 566782 494041 566842 494101
rect 566902 494041 566962 494101
rect 567022 494041 567082 494101
rect 567142 494041 567202 494101
rect 567262 494041 567322 494101
rect 567382 494041 567442 494101
rect 567502 494041 567562 494101
rect 572332 494176 572392 494236
rect 572452 494176 572512 494236
rect 572572 494176 572632 494236
rect 572692 494176 572752 494236
rect 572812 494176 572872 494236
rect 572932 494176 572992 494236
rect 573052 494176 573112 494236
rect 573172 494176 573232 494236
rect 573292 494176 573352 494236
rect 573412 494176 573472 494236
rect 573532 494176 573592 494236
rect 573652 494176 573712 494236
rect 573772 494176 573832 494236
rect 573892 494176 573952 494236
rect 574012 494176 574072 494236
rect 574132 494176 574192 494236
rect 574252 494176 574312 494236
rect 574372 494176 574432 494236
rect 574492 494176 574552 494236
rect 574612 494176 574672 494236
rect 574732 494176 574792 494236
rect 574852 494176 574912 494236
rect 574972 494176 575032 494236
rect 575092 494176 575152 494236
rect 575212 494176 575272 494236
rect 575332 494176 575392 494236
rect 575452 494176 575512 494236
rect 575572 494176 575632 494236
rect 575692 494176 575752 494236
rect 575812 494176 575872 494236
rect 575932 494176 575992 494236
rect 576052 494176 576112 494236
rect 576172 494176 576232 494236
rect 576292 494176 576352 494236
rect 576412 494176 576472 494236
rect 576532 494176 576592 494236
rect 576652 494176 576712 494236
rect 576772 494176 576832 494236
rect 576892 494176 576952 494236
rect 577012 494176 577072 494236
rect 577132 494176 577192 494236
rect 577252 494176 577312 494236
rect 577372 494176 577432 494236
rect 577492 494176 577552 494236
rect 577612 494176 577672 494236
rect 572332 494056 572392 494116
rect 572452 494056 572512 494116
rect 572572 494056 572632 494116
rect 572692 494056 572752 494116
rect 572812 494056 572872 494116
rect 572932 494056 572992 494116
rect 573052 494056 573112 494116
rect 573172 494056 573232 494116
rect 573292 494056 573352 494116
rect 573412 494056 573472 494116
rect 573532 494056 573592 494116
rect 573652 494056 573712 494116
rect 573772 494056 573832 494116
rect 573892 494056 573952 494116
rect 574012 494056 574072 494116
rect 574132 494056 574192 494116
rect 574252 494056 574312 494116
rect 574372 494056 574432 494116
rect 574492 494056 574552 494116
rect 574612 494056 574672 494116
rect 574732 494056 574792 494116
rect 574852 494056 574912 494116
rect 574972 494056 575032 494116
rect 575092 494056 575152 494116
rect 575212 494056 575272 494116
rect 575332 494056 575392 494116
rect 575452 494056 575512 494116
rect 575572 494056 575632 494116
rect 575692 494056 575752 494116
rect 575812 494056 575872 494116
rect 575932 494056 575992 494116
rect 576052 494056 576112 494116
rect 576172 494056 576232 494116
rect 576292 494056 576352 494116
rect 576412 494056 576472 494116
rect 576532 494056 576592 494116
rect 576652 494056 576712 494116
rect 576772 494056 576832 494116
rect 576892 494056 576952 494116
rect 577012 494056 577072 494116
rect 577132 494056 577192 494116
rect 577252 494056 577312 494116
rect 577372 494056 577432 494116
rect 577492 494056 577552 494116
rect 577612 494056 577672 494116
rect 503920 475206 504020 475306
rect 504144 475206 504244 475306
rect 504368 475206 504468 475306
rect 504592 475206 504692 475306
rect 504816 475206 504916 475306
rect 505040 475206 505140 475306
rect 505264 475206 505364 475306
rect 505488 475206 505588 475306
rect 505712 475206 505812 475306
rect 505936 475206 506036 475306
rect 506160 475206 506260 475306
rect 506384 475206 506484 475306
rect 506608 475206 506708 475306
rect 506832 475206 506932 475306
rect 507056 475206 507156 475306
rect 507280 475206 507380 475306
rect 507504 475206 507604 475306
rect 507728 475206 507828 475306
rect 507952 475206 508052 475306
rect 508176 475206 508276 475306
rect 508400 475206 508500 475306
rect 508624 475206 508724 475306
rect 508848 475206 508948 475306
rect 509072 475206 509172 475306
rect 509296 475206 509396 475306
rect 509520 475206 509620 475306
rect 509744 475206 509844 475306
rect 509968 475206 510068 475306
rect 510192 475206 510292 475306
rect 510416 475206 510516 475306
rect 503920 474982 504020 475082
rect 504144 474982 504244 475082
rect 504368 474982 504468 475082
rect 504592 474982 504692 475082
rect 504816 474982 504916 475082
rect 505040 474982 505140 475082
rect 505264 474982 505364 475082
rect 505488 474982 505588 475082
rect 505712 474982 505812 475082
rect 505936 474982 506036 475082
rect 506160 474982 506260 475082
rect 506384 474982 506484 475082
rect 506608 474982 506708 475082
rect 506832 474982 506932 475082
rect 507056 474982 507156 475082
rect 507280 474982 507380 475082
rect 507504 474982 507604 475082
rect 507728 474982 507828 475082
rect 507952 474982 508052 475082
rect 508176 474982 508276 475082
rect 508400 474982 508500 475082
rect 508624 474982 508724 475082
rect 508848 474982 508948 475082
rect 509072 474982 509172 475082
rect 509296 474982 509396 475082
rect 509520 474982 509620 475082
rect 509744 474982 509844 475082
rect 509968 474982 510068 475082
rect 510192 474982 510292 475082
rect 510416 474982 510516 475082
rect 503920 474758 504020 474858
rect 504144 474758 504244 474858
rect 504368 474758 504468 474858
rect 504592 474758 504692 474858
rect 504816 474758 504916 474858
rect 505040 474758 505140 474858
rect 505264 474758 505364 474858
rect 505488 474758 505588 474858
rect 505712 474758 505812 474858
rect 505936 474758 506036 474858
rect 506160 474758 506260 474858
rect 506384 474758 506484 474858
rect 506608 474758 506708 474858
rect 506832 474758 506932 474858
rect 507056 474758 507156 474858
rect 507280 474758 507380 474858
rect 507504 474758 507604 474858
rect 507728 474758 507828 474858
rect 507952 474758 508052 474858
rect 508176 474758 508276 474858
rect 508400 474758 508500 474858
rect 508624 474758 508724 474858
rect 508848 474758 508948 474858
rect 509072 474758 509172 474858
rect 509296 474758 509396 474858
rect 509520 474758 509620 474858
rect 509744 474758 509844 474858
rect 509968 474758 510068 474858
rect 510192 474758 510292 474858
rect 510416 474758 510516 474858
rect 503920 474534 504020 474634
rect 504144 474534 504244 474634
rect 504368 474534 504468 474634
rect 504592 474534 504692 474634
rect 504816 474534 504916 474634
rect 505040 474534 505140 474634
rect 505264 474534 505364 474634
rect 505488 474534 505588 474634
rect 505712 474534 505812 474634
rect 505936 474534 506036 474634
rect 506160 474534 506260 474634
rect 506384 474534 506484 474634
rect 506608 474534 506708 474634
rect 506832 474534 506932 474634
rect 507056 474534 507156 474634
rect 507280 474534 507380 474634
rect 507504 474534 507604 474634
rect 507728 474534 507828 474634
rect 507952 474534 508052 474634
rect 508176 474534 508276 474634
rect 508400 474534 508500 474634
rect 508624 474534 508724 474634
rect 508848 474534 508948 474634
rect 509072 474534 509172 474634
rect 509296 474534 509396 474634
rect 509520 474534 509620 474634
rect 509744 474534 509844 474634
rect 509968 474534 510068 474634
rect 510192 474534 510292 474634
rect 510416 474534 510516 474634
rect 500398 474180 500498 474280
rect 500622 474180 500722 474280
rect 500846 474180 500946 474280
rect 501070 474180 501170 474280
rect 501294 474180 501394 474280
rect 503920 474310 504020 474410
rect 504144 474310 504244 474410
rect 504368 474310 504468 474410
rect 504592 474310 504692 474410
rect 504816 474310 504916 474410
rect 505040 474310 505140 474410
rect 505264 474310 505364 474410
rect 505488 474310 505588 474410
rect 505712 474310 505812 474410
rect 505936 474310 506036 474410
rect 506160 474310 506260 474410
rect 506384 474310 506484 474410
rect 506608 474310 506708 474410
rect 506832 474310 506932 474410
rect 507056 474310 507156 474410
rect 507280 474310 507380 474410
rect 507504 474310 507604 474410
rect 507728 474310 507828 474410
rect 507952 474310 508052 474410
rect 508176 474310 508276 474410
rect 508400 474310 508500 474410
rect 508624 474310 508724 474410
rect 508848 474310 508948 474410
rect 509072 474310 509172 474410
rect 509296 474310 509396 474410
rect 509520 474310 509620 474410
rect 509744 474310 509844 474410
rect 509968 474310 510068 474410
rect 510192 474310 510292 474410
rect 510416 474310 510516 474410
rect 517320 475206 517420 475306
rect 517544 475206 517644 475306
rect 517768 475206 517868 475306
rect 517992 475206 518092 475306
rect 518216 475206 518316 475306
rect 518440 475206 518540 475306
rect 518664 475206 518764 475306
rect 518888 475206 518988 475306
rect 519112 475206 519212 475306
rect 519336 475206 519436 475306
rect 519560 475206 519660 475306
rect 519784 475206 519884 475306
rect 520008 475206 520108 475306
rect 520232 475206 520332 475306
rect 520456 475206 520556 475306
rect 520680 475206 520780 475306
rect 520904 475206 521004 475306
rect 521128 475206 521228 475306
rect 521352 475206 521452 475306
rect 521576 475206 521676 475306
rect 521800 475206 521900 475306
rect 522024 475206 522124 475306
rect 522248 475206 522348 475306
rect 522472 475206 522572 475306
rect 522696 475206 522796 475306
rect 522920 475206 523020 475306
rect 523144 475206 523244 475306
rect 523368 475206 523468 475306
rect 523592 475206 523692 475306
rect 523816 475206 523916 475306
rect 517320 474982 517420 475082
rect 517544 474982 517644 475082
rect 517768 474982 517868 475082
rect 517992 474982 518092 475082
rect 518216 474982 518316 475082
rect 518440 474982 518540 475082
rect 518664 474982 518764 475082
rect 518888 474982 518988 475082
rect 519112 474982 519212 475082
rect 519336 474982 519436 475082
rect 519560 474982 519660 475082
rect 519784 474982 519884 475082
rect 520008 474982 520108 475082
rect 520232 474982 520332 475082
rect 520456 474982 520556 475082
rect 520680 474982 520780 475082
rect 520904 474982 521004 475082
rect 521128 474982 521228 475082
rect 521352 474982 521452 475082
rect 521576 474982 521676 475082
rect 521800 474982 521900 475082
rect 522024 474982 522124 475082
rect 522248 474982 522348 475082
rect 522472 474982 522572 475082
rect 522696 474982 522796 475082
rect 522920 474982 523020 475082
rect 523144 474982 523244 475082
rect 523368 474982 523468 475082
rect 523592 474982 523692 475082
rect 523816 474982 523916 475082
rect 517320 474758 517420 474858
rect 517544 474758 517644 474858
rect 517768 474758 517868 474858
rect 517992 474758 518092 474858
rect 518216 474758 518316 474858
rect 518440 474758 518540 474858
rect 518664 474758 518764 474858
rect 518888 474758 518988 474858
rect 519112 474758 519212 474858
rect 519336 474758 519436 474858
rect 519560 474758 519660 474858
rect 519784 474758 519884 474858
rect 520008 474758 520108 474858
rect 520232 474758 520332 474858
rect 520456 474758 520556 474858
rect 520680 474758 520780 474858
rect 520904 474758 521004 474858
rect 521128 474758 521228 474858
rect 521352 474758 521452 474858
rect 521576 474758 521676 474858
rect 521800 474758 521900 474858
rect 522024 474758 522124 474858
rect 522248 474758 522348 474858
rect 522472 474758 522572 474858
rect 522696 474758 522796 474858
rect 522920 474758 523020 474858
rect 523144 474758 523244 474858
rect 523368 474758 523468 474858
rect 523592 474758 523692 474858
rect 523816 474758 523916 474858
rect 517320 474534 517420 474634
rect 517544 474534 517644 474634
rect 517768 474534 517868 474634
rect 517992 474534 518092 474634
rect 518216 474534 518316 474634
rect 518440 474534 518540 474634
rect 518664 474534 518764 474634
rect 518888 474534 518988 474634
rect 519112 474534 519212 474634
rect 519336 474534 519436 474634
rect 519560 474534 519660 474634
rect 519784 474534 519884 474634
rect 520008 474534 520108 474634
rect 520232 474534 520332 474634
rect 520456 474534 520556 474634
rect 520680 474534 520780 474634
rect 520904 474534 521004 474634
rect 521128 474534 521228 474634
rect 521352 474534 521452 474634
rect 521576 474534 521676 474634
rect 521800 474534 521900 474634
rect 522024 474534 522124 474634
rect 522248 474534 522348 474634
rect 522472 474534 522572 474634
rect 522696 474534 522796 474634
rect 522920 474534 523020 474634
rect 523144 474534 523244 474634
rect 523368 474534 523468 474634
rect 523592 474534 523692 474634
rect 523816 474534 523916 474634
rect 517320 474310 517420 474410
rect 517544 474310 517644 474410
rect 517768 474310 517868 474410
rect 517992 474310 518092 474410
rect 518216 474310 518316 474410
rect 518440 474310 518540 474410
rect 518664 474310 518764 474410
rect 518888 474310 518988 474410
rect 519112 474310 519212 474410
rect 519336 474310 519436 474410
rect 519560 474310 519660 474410
rect 519784 474310 519884 474410
rect 520008 474310 520108 474410
rect 520232 474310 520332 474410
rect 520456 474310 520556 474410
rect 520680 474310 520780 474410
rect 520904 474310 521004 474410
rect 521128 474310 521228 474410
rect 521352 474310 521452 474410
rect 521576 474310 521676 474410
rect 521800 474310 521900 474410
rect 522024 474310 522124 474410
rect 522248 474310 522348 474410
rect 522472 474310 522572 474410
rect 522696 474310 522796 474410
rect 522920 474310 523020 474410
rect 523144 474310 523244 474410
rect 523368 474310 523468 474410
rect 523592 474310 523692 474410
rect 523816 474310 523916 474410
rect 500398 473956 500498 474056
rect 500622 473956 500722 474056
rect 500846 473956 500946 474056
rect 501070 473956 501170 474056
rect 501294 473956 501394 474056
rect 500398 473732 500498 473832
rect 500622 473732 500722 473832
rect 500846 473732 500946 473832
rect 501070 473732 501170 473832
rect 501294 473732 501394 473832
rect 500398 473508 500498 473608
rect 500622 473508 500722 473608
rect 500846 473508 500946 473608
rect 501070 473508 501170 473608
rect 501294 473508 501394 473608
rect 500398 473284 500498 473384
rect 500622 473284 500722 473384
rect 500846 473284 500946 473384
rect 501070 473284 501170 473384
rect 501294 473284 501394 473384
rect 500398 473060 500498 473160
rect 500622 473060 500722 473160
rect 500846 473060 500946 473160
rect 501070 473060 501170 473160
rect 501294 473060 501394 473160
rect 500398 472836 500498 472936
rect 500622 472836 500722 472936
rect 500846 472836 500946 472936
rect 501070 472836 501170 472936
rect 501294 472836 501394 472936
rect 500398 472612 500498 472712
rect 500622 472612 500722 472712
rect 500846 472612 500946 472712
rect 501070 472612 501170 472712
rect 501294 472612 501394 472712
rect 527618 474180 527718 474280
rect 527842 474180 527942 474280
rect 528066 474180 528166 474280
rect 528290 474180 528390 474280
rect 528514 474180 528614 474280
rect 527618 473956 527718 474056
rect 527842 473956 527942 474056
rect 528066 473956 528166 474056
rect 528290 473956 528390 474056
rect 528514 473956 528614 474056
rect 527618 473732 527718 473832
rect 527842 473732 527942 473832
rect 528066 473732 528166 473832
rect 528290 473732 528390 473832
rect 528514 473732 528614 473832
rect 527618 473508 527718 473608
rect 527842 473508 527942 473608
rect 528066 473508 528166 473608
rect 528290 473508 528390 473608
rect 528514 473508 528614 473608
rect 527618 473284 527718 473384
rect 527842 473284 527942 473384
rect 528066 473284 528166 473384
rect 528290 473284 528390 473384
rect 528514 473284 528614 473384
rect 527618 473060 527718 473160
rect 527842 473060 527942 473160
rect 528066 473060 528166 473160
rect 528290 473060 528390 473160
rect 528514 473060 528614 473160
rect 527618 472836 527718 472936
rect 527842 472836 527942 472936
rect 528066 472836 528166 472936
rect 528290 472836 528390 472936
rect 528514 472836 528614 472936
rect 527618 472612 527718 472712
rect 527842 472612 527942 472712
rect 528066 472612 528166 472712
rect 528290 472612 528390 472712
rect 528514 472612 528614 472712
rect 500398 472388 500498 472488
rect 500622 472388 500722 472488
rect 500846 472388 500946 472488
rect 501070 472388 501170 472488
rect 501294 472388 501394 472488
rect 500398 472164 500498 472264
rect 500622 472164 500722 472264
rect 500846 472164 500946 472264
rect 501070 472164 501170 472264
rect 501294 472164 501394 472264
rect 500398 471940 500498 472040
rect 500622 471940 500722 472040
rect 500846 471940 500946 472040
rect 501070 471940 501170 472040
rect 501294 471940 501394 472040
rect 500398 471716 500498 471816
rect 500622 471716 500722 471816
rect 500846 471716 500946 471816
rect 501070 471716 501170 471816
rect 501294 471716 501394 471816
rect 500398 471492 500498 471592
rect 500622 471492 500722 471592
rect 500846 471492 500946 471592
rect 501070 471492 501170 471592
rect 501294 471492 501394 471592
rect 500398 471268 500498 471368
rect 500622 471268 500722 471368
rect 500846 471268 500946 471368
rect 501070 471268 501170 471368
rect 501294 471268 501394 471368
rect 500398 471044 500498 471144
rect 500622 471044 500722 471144
rect 500846 471044 500946 471144
rect 501070 471044 501170 471144
rect 501294 471044 501394 471144
rect 500398 470820 500498 470920
rect 500622 470820 500722 470920
rect 500846 470820 500946 470920
rect 501070 470820 501170 470920
rect 501294 470820 501394 470920
rect 500398 470596 500498 470696
rect 500622 470596 500722 470696
rect 500846 470596 500946 470696
rect 501070 470596 501170 470696
rect 501294 470596 501394 470696
rect 500398 470372 500498 470472
rect 500622 470372 500722 470472
rect 500846 470372 500946 470472
rect 501070 470372 501170 470472
rect 501294 470372 501394 470472
rect 500398 470148 500498 470248
rect 500622 470148 500722 470248
rect 500846 470148 500946 470248
rect 501070 470148 501170 470248
rect 501294 470148 501394 470248
rect 500398 469924 500498 470024
rect 500622 469924 500722 470024
rect 500846 469924 500946 470024
rect 501070 469924 501170 470024
rect 501294 469924 501394 470024
rect 500398 469700 500498 469800
rect 500622 469700 500722 469800
rect 500846 469700 500946 469800
rect 501070 469700 501170 469800
rect 501294 469700 501394 469800
rect 500398 469476 500498 469576
rect 500622 469476 500722 469576
rect 500846 469476 500946 469576
rect 501070 469476 501170 469576
rect 501294 469476 501394 469576
rect 500398 469252 500498 469352
rect 500622 469252 500722 469352
rect 500846 469252 500946 469352
rect 501070 469252 501170 469352
rect 501294 469252 501394 469352
rect 500398 469028 500498 469128
rect 500622 469028 500722 469128
rect 500846 469028 500946 469128
rect 501070 469028 501170 469128
rect 501294 469028 501394 469128
rect 500398 468804 500498 468904
rect 500622 468804 500722 468904
rect 500846 468804 500946 468904
rect 501070 468804 501170 468904
rect 501294 468804 501394 468904
rect 500398 468580 500498 468680
rect 500622 468580 500722 468680
rect 500846 468580 500946 468680
rect 501070 468580 501170 468680
rect 501294 468580 501394 468680
rect 500398 468356 500498 468456
rect 500622 468356 500722 468456
rect 500846 468356 500946 468456
rect 501070 468356 501170 468456
rect 501294 468356 501394 468456
rect 500398 468132 500498 468232
rect 500622 468132 500722 468232
rect 500846 468132 500946 468232
rect 501070 468132 501170 468232
rect 501294 468132 501394 468232
rect 500398 467908 500498 468008
rect 500622 467908 500722 468008
rect 500846 467908 500946 468008
rect 501070 467908 501170 468008
rect 501294 467908 501394 468008
rect 500398 467684 500498 467784
rect 500622 467684 500722 467784
rect 500846 467684 500946 467784
rect 501070 467684 501170 467784
rect 501294 467684 501394 467784
rect 500398 463710 500498 463810
rect 500622 463710 500722 463810
rect 500846 463710 500946 463810
rect 501070 463710 501170 463810
rect 501294 463710 501394 463810
rect 500398 463486 500498 463586
rect 500622 463486 500722 463586
rect 500846 463486 500946 463586
rect 501070 463486 501170 463586
rect 501294 463486 501394 463586
rect 500398 463262 500498 463362
rect 500622 463262 500722 463362
rect 500846 463262 500946 463362
rect 501070 463262 501170 463362
rect 501294 463262 501394 463362
rect 500398 463038 500498 463138
rect 500622 463038 500722 463138
rect 500846 463038 500946 463138
rect 501070 463038 501170 463138
rect 501294 463038 501394 463138
rect 500398 462814 500498 462914
rect 500622 462814 500722 462914
rect 500846 462814 500946 462914
rect 501070 462814 501170 462914
rect 501294 462814 501394 462914
rect 500398 462590 500498 462690
rect 500622 462590 500722 462690
rect 500846 462590 500946 462690
rect 501070 462590 501170 462690
rect 501294 462590 501394 462690
rect 500398 462366 500498 462466
rect 500622 462366 500722 462466
rect 500846 462366 500946 462466
rect 501070 462366 501170 462466
rect 501294 462366 501394 462466
rect 500398 462142 500498 462242
rect 500622 462142 500722 462242
rect 500846 462142 500946 462242
rect 501070 462142 501170 462242
rect 501294 462142 501394 462242
rect 500398 461918 500498 462018
rect 500622 461918 500722 462018
rect 500846 461918 500946 462018
rect 501070 461918 501170 462018
rect 501294 461918 501394 462018
rect 500398 461694 500498 461794
rect 500622 461694 500722 461794
rect 500846 461694 500946 461794
rect 501070 461694 501170 461794
rect 501294 461694 501394 461794
rect 500398 461470 500498 461570
rect 500622 461470 500722 461570
rect 500846 461470 500946 461570
rect 501070 461470 501170 461570
rect 501294 461470 501394 461570
rect 500398 461246 500498 461346
rect 500622 461246 500722 461346
rect 500846 461246 500946 461346
rect 501070 461246 501170 461346
rect 501294 461246 501394 461346
rect 500398 461022 500498 461122
rect 500622 461022 500722 461122
rect 500846 461022 500946 461122
rect 501070 461022 501170 461122
rect 501294 461022 501394 461122
rect 502868 470192 502982 470210
rect 502868 470140 502874 470192
rect 502874 470140 502978 470192
rect 502978 470140 502982 470192
rect 502868 469570 502982 470140
rect 502868 469518 502874 469570
rect 502874 469518 502978 469570
rect 502978 469518 502982 469570
rect 502868 469112 502982 469518
rect 502868 469060 502874 469112
rect 502874 469060 502978 469112
rect 502978 469060 502982 469112
rect 502868 468536 502982 469060
rect 502868 468484 502874 468536
rect 502874 468484 502978 468536
rect 502978 468484 502982 468536
rect 502868 467964 502982 468484
rect 502868 467912 502874 467964
rect 502874 467912 502978 467964
rect 502978 467912 502982 467964
rect 502868 467392 502982 467912
rect 502868 467340 502874 467392
rect 502874 467340 502978 467392
rect 502978 467340 502982 467392
rect 502868 466820 502982 467340
rect 502868 466768 502874 466820
rect 502874 466768 502978 466820
rect 502978 466768 502982 466820
rect 502868 466248 502982 466768
rect 502868 466196 502874 466248
rect 502874 466196 502978 466248
rect 502978 466196 502982 466248
rect 502868 465676 502982 466196
rect 502868 465624 502874 465676
rect 502874 465624 502978 465676
rect 502978 465624 502982 465676
rect 502868 465104 502982 465624
rect 502868 465052 502874 465104
rect 502874 465052 502978 465104
rect 502978 465052 502982 465104
rect 502868 464532 502982 465052
rect 502868 464480 502874 464532
rect 502874 464480 502978 464532
rect 502978 464480 502982 464532
rect 502868 463960 502982 464480
rect 502868 463908 502874 463960
rect 502874 463908 502978 463960
rect 502978 463908 502982 463960
rect 502868 463388 502982 463908
rect 502868 463336 502874 463388
rect 502874 463336 502978 463388
rect 502978 463336 502982 463388
rect 502868 462816 502982 463336
rect 502868 462764 502874 462816
rect 502874 462764 502978 462816
rect 502978 462764 502982 462816
rect 502868 462244 502982 462764
rect 502868 462192 502874 462244
rect 502874 462192 502978 462244
rect 502978 462192 502982 462244
rect 502868 462134 502982 462192
rect 502868 462082 502874 462134
rect 502874 462082 502978 462134
rect 502978 462082 502982 462134
rect 502868 461676 502982 462082
rect 502868 461624 502874 461676
rect 502874 461624 502978 461676
rect 502978 461624 502982 461676
rect 502868 461064 502982 461624
rect 502868 461012 502874 461064
rect 502874 461012 502978 461064
rect 502978 461012 502982 461064
rect 502868 460964 502982 461012
rect 505803 468952 506055 469552
rect 511770 470116 511830 470176
rect 511890 470116 511950 470176
rect 511770 469996 511830 470056
rect 511890 469996 511950 470056
rect 511770 469876 511830 469936
rect 511890 469876 511950 469936
rect 511770 469756 511830 469816
rect 511890 469756 511950 469816
rect 511770 469636 511830 469696
rect 511890 469636 511950 469696
rect 500398 460798 500498 460898
rect 500622 460798 500722 460898
rect 500846 460798 500946 460898
rect 501070 460798 501170 460898
rect 501294 460798 501394 460898
rect 500398 460574 500498 460674
rect 500622 460574 500722 460674
rect 500846 460574 500946 460674
rect 501070 460574 501170 460674
rect 501294 460574 501394 460674
rect 505803 460461 506055 461061
rect 525660 472498 526498 472504
rect 525660 461254 525666 472498
rect 525666 461254 526492 472498
rect 526492 461254 526498 472498
rect 525660 461248 526498 461254
rect 527618 472388 527718 472488
rect 527842 472388 527942 472488
rect 528066 472388 528166 472488
rect 528290 472388 528390 472488
rect 528514 472388 528614 472488
rect 527618 472164 527718 472264
rect 527842 472164 527942 472264
rect 528066 472164 528166 472264
rect 528290 472164 528390 472264
rect 528514 472164 528614 472264
rect 527618 471940 527718 472040
rect 527842 471940 527942 472040
rect 528066 471940 528166 472040
rect 528290 471940 528390 472040
rect 528514 471940 528614 472040
rect 527618 471716 527718 471816
rect 527842 471716 527942 471816
rect 528066 471716 528166 471816
rect 528290 471716 528390 471816
rect 528514 471716 528614 471816
rect 527618 471492 527718 471592
rect 527842 471492 527942 471592
rect 528066 471492 528166 471592
rect 528290 471492 528390 471592
rect 528514 471492 528614 471592
rect 527618 471268 527718 471368
rect 527842 471268 527942 471368
rect 528066 471268 528166 471368
rect 528290 471268 528390 471368
rect 528514 471268 528614 471368
rect 527618 471044 527718 471144
rect 527842 471044 527942 471144
rect 528066 471044 528166 471144
rect 528290 471044 528390 471144
rect 528514 471044 528614 471144
rect 527618 470820 527718 470920
rect 527842 470820 527942 470920
rect 528066 470820 528166 470920
rect 528290 470820 528390 470920
rect 528514 470820 528614 470920
rect 527618 470596 527718 470696
rect 527842 470596 527942 470696
rect 528066 470596 528166 470696
rect 528290 470596 528390 470696
rect 528514 470596 528614 470696
rect 527618 470372 527718 470472
rect 527842 470372 527942 470472
rect 528066 470372 528166 470472
rect 528290 470372 528390 470472
rect 528514 470372 528614 470472
rect 527618 470148 527718 470248
rect 527842 470148 527942 470248
rect 528066 470148 528166 470248
rect 528290 470148 528390 470248
rect 528514 470148 528614 470248
rect 527618 469924 527718 470024
rect 527842 469924 527942 470024
rect 528066 469924 528166 470024
rect 528290 469924 528390 470024
rect 528514 469924 528614 470024
rect 527618 469700 527718 469800
rect 527842 469700 527942 469800
rect 528066 469700 528166 469800
rect 528290 469700 528390 469800
rect 528514 469700 528614 469800
rect 527618 469476 527718 469576
rect 527842 469476 527942 469576
rect 528066 469476 528166 469576
rect 528290 469476 528390 469576
rect 528514 469476 528614 469576
rect 527618 469252 527718 469352
rect 527842 469252 527942 469352
rect 528066 469252 528166 469352
rect 528290 469252 528390 469352
rect 528514 469252 528614 469352
rect 527618 469028 527718 469128
rect 527842 469028 527942 469128
rect 528066 469028 528166 469128
rect 528290 469028 528390 469128
rect 528514 469028 528614 469128
rect 527618 468804 527718 468904
rect 527842 468804 527942 468904
rect 528066 468804 528166 468904
rect 528290 468804 528390 468904
rect 528514 468804 528614 468904
rect 527618 468580 527718 468680
rect 527842 468580 527942 468680
rect 528066 468580 528166 468680
rect 528290 468580 528390 468680
rect 528514 468580 528614 468680
rect 527618 468356 527718 468456
rect 527842 468356 527942 468456
rect 528066 468356 528166 468456
rect 528290 468356 528390 468456
rect 528514 468356 528614 468456
rect 527618 468132 527718 468232
rect 527842 468132 527942 468232
rect 528066 468132 528166 468232
rect 528290 468132 528390 468232
rect 528514 468132 528614 468232
rect 527618 467908 527718 468008
rect 527842 467908 527942 468008
rect 528066 467908 528166 468008
rect 528290 467908 528390 468008
rect 528514 467908 528614 468008
rect 527618 467684 527718 467784
rect 527842 467684 527942 467784
rect 528066 467684 528166 467784
rect 528290 467684 528390 467784
rect 528514 467684 528614 467784
rect 527618 463710 527718 463810
rect 527842 463710 527942 463810
rect 528066 463710 528166 463810
rect 528290 463710 528390 463810
rect 528514 463710 528614 463810
rect 527618 463486 527718 463586
rect 527842 463486 527942 463586
rect 528066 463486 528166 463586
rect 528290 463486 528390 463586
rect 528514 463486 528614 463586
rect 527618 463262 527718 463362
rect 527842 463262 527942 463362
rect 528066 463262 528166 463362
rect 528290 463262 528390 463362
rect 528514 463262 528614 463362
rect 527618 463038 527718 463138
rect 527842 463038 527942 463138
rect 528066 463038 528166 463138
rect 528290 463038 528390 463138
rect 528514 463038 528614 463138
rect 527618 462814 527718 462914
rect 527842 462814 527942 462914
rect 528066 462814 528166 462914
rect 528290 462814 528390 462914
rect 528514 462814 528614 462914
rect 527618 462590 527718 462690
rect 527842 462590 527942 462690
rect 528066 462590 528166 462690
rect 528290 462590 528390 462690
rect 528514 462590 528614 462690
rect 527618 462366 527718 462466
rect 527842 462366 527942 462466
rect 528066 462366 528166 462466
rect 528290 462366 528390 462466
rect 528514 462366 528614 462466
rect 527618 462142 527718 462242
rect 527842 462142 527942 462242
rect 528066 462142 528166 462242
rect 528290 462142 528390 462242
rect 528514 462142 528614 462242
rect 527618 461918 527718 462018
rect 527842 461918 527942 462018
rect 528066 461918 528166 462018
rect 528290 461918 528390 462018
rect 528514 461918 528614 462018
rect 527618 461694 527718 461794
rect 527842 461694 527942 461794
rect 528066 461694 528166 461794
rect 528290 461694 528390 461794
rect 528514 461694 528614 461794
rect 527618 461470 527718 461570
rect 527842 461470 527942 461570
rect 528066 461470 528166 461570
rect 528290 461470 528390 461570
rect 528514 461470 528614 461570
rect 527618 461246 527718 461346
rect 527842 461246 527942 461346
rect 528066 461246 528166 461346
rect 528290 461246 528390 461346
rect 528514 461246 528614 461346
rect 500398 460350 500498 460450
rect 500622 460350 500722 460450
rect 500846 460350 500946 460450
rect 501070 460350 501170 460450
rect 501294 460350 501394 460450
rect 500398 460126 500498 460226
rect 500622 460126 500722 460226
rect 500846 460126 500946 460226
rect 501070 460126 501170 460226
rect 501294 460126 501394 460226
rect 500398 459902 500498 460002
rect 500622 459902 500722 460002
rect 500846 459902 500946 460002
rect 501070 459902 501170 460002
rect 501294 459902 501394 460002
rect 500398 459678 500498 459778
rect 500622 459678 500722 459778
rect 500846 459678 500946 459778
rect 501070 459678 501170 459778
rect 501294 459678 501394 459778
rect 500398 459454 500498 459554
rect 500622 459454 500722 459554
rect 500846 459454 500946 459554
rect 501070 459454 501170 459554
rect 501294 459454 501394 459554
rect 500398 459230 500498 459330
rect 500622 459230 500722 459330
rect 500846 459230 500946 459330
rect 501070 459230 501170 459330
rect 501294 459230 501394 459330
rect 500398 459006 500498 459106
rect 500622 459006 500722 459106
rect 500846 459006 500946 459106
rect 501070 459006 501170 459106
rect 501294 459006 501394 459106
rect 500398 458782 500498 458882
rect 500622 458782 500722 458882
rect 500846 458782 500946 458882
rect 501070 458782 501170 458882
rect 501294 458782 501394 458882
rect 500398 458558 500498 458658
rect 500622 458558 500722 458658
rect 500846 458558 500946 458658
rect 501070 458558 501170 458658
rect 501294 458558 501394 458658
rect 500398 458334 500498 458434
rect 500622 458334 500722 458434
rect 500846 458334 500946 458434
rect 501070 458334 501170 458434
rect 501294 458334 501394 458434
rect 500398 458110 500498 458210
rect 500622 458110 500722 458210
rect 500846 458110 500946 458210
rect 501070 458110 501170 458210
rect 501294 458110 501394 458210
rect 500398 457886 500498 457986
rect 500622 457886 500722 457986
rect 500846 457886 500946 457986
rect 501070 457886 501170 457986
rect 501294 457886 501394 457986
rect 500398 457662 500498 457762
rect 500622 457662 500722 457762
rect 500846 457662 500946 457762
rect 501070 457662 501170 457762
rect 501294 457662 501394 457762
rect 500398 457438 500498 457538
rect 500622 457438 500722 457538
rect 500846 457438 500946 457538
rect 501070 457438 501170 457538
rect 501294 457438 501394 457538
rect 500398 457214 500498 457314
rect 500622 457214 500722 457314
rect 500846 457214 500946 457314
rect 501070 457214 501170 457314
rect 501294 457214 501394 457314
rect 502432 460352 502750 460446
rect 502432 459952 502528 460352
rect 502528 459952 502628 460352
rect 502628 459952 502750 460352
rect 502432 458862 502750 459952
rect 502432 458782 502668 458862
rect 502668 458782 502748 458862
rect 502748 458782 502750 458862
rect 502432 457942 502750 458782
rect 502432 457862 502668 457942
rect 502668 457862 502748 457942
rect 502748 457862 502750 457942
rect 502432 457022 502750 457862
rect 502432 456942 502668 457022
rect 502668 456942 502748 457022
rect 502748 456942 502750 457022
rect 502432 456102 502750 456942
rect 502432 456022 502668 456102
rect 502668 456022 502748 456102
rect 502748 456022 502750 456102
rect 502432 455182 502750 456022
rect 502432 455102 502668 455182
rect 502668 455102 502748 455182
rect 502748 455102 502750 455182
rect 502432 454442 502750 455102
rect 502432 454042 502528 454442
rect 502528 454042 502628 454442
rect 502628 454042 502750 454442
rect 502432 453362 502750 454042
rect 502432 453282 502668 453362
rect 502668 453282 502748 453362
rect 502748 453282 502750 453362
rect 502432 452442 502750 453282
rect 502432 452362 502668 452442
rect 502668 452362 502748 452442
rect 502748 452362 502750 452442
rect 502432 451522 502750 452362
rect 502432 451442 502668 451522
rect 502668 451442 502748 451522
rect 502748 451442 502750 451522
rect 502432 450602 502750 451442
rect 502432 450522 502668 450602
rect 502668 450522 502748 450602
rect 502748 450522 502750 450602
rect 502432 449682 502750 450522
rect 502432 449602 502668 449682
rect 502668 449602 502748 449682
rect 502748 449602 502750 449682
rect 502432 448942 502750 449602
rect 502432 448542 502528 448942
rect 502528 448542 502628 448942
rect 502628 448542 502750 448942
rect 502432 447862 502750 448542
rect 502432 447782 502668 447862
rect 502668 447782 502748 447862
rect 502748 447782 502750 447862
rect 502432 446942 502750 447782
rect 502432 446862 502668 446942
rect 502668 446862 502748 446942
rect 502748 446862 502750 446942
rect 502432 446022 502750 446862
rect 502432 445942 502668 446022
rect 502668 445942 502748 446022
rect 502748 445942 502750 446022
rect 502432 445102 502750 445942
rect 502432 445022 502668 445102
rect 502668 445022 502748 445102
rect 502748 445022 502750 445102
rect 502432 444182 502750 445022
rect 502432 444102 502668 444182
rect 502668 444102 502748 444182
rect 502748 444102 502750 444182
rect 502432 442986 502750 444102
rect 502432 442586 502526 442986
rect 502526 442586 502626 442986
rect 502626 442586 502750 442986
rect 502432 442508 502750 442586
rect 527618 461022 527718 461122
rect 527842 461022 527942 461122
rect 528066 461022 528166 461122
rect 528290 461022 528390 461122
rect 528514 461022 528614 461122
rect 500418 437440 500518 437540
rect 500642 437440 500742 437540
rect 500866 437440 500966 437540
rect 501090 437440 501190 437540
rect 501314 437440 501414 437540
rect 500418 437216 500518 437316
rect 500642 437216 500742 437316
rect 500866 437216 500966 437316
rect 501090 437216 501190 437316
rect 501314 437216 501414 437316
rect 500418 436992 500518 437092
rect 500642 436992 500742 437092
rect 500866 436992 500966 437092
rect 501090 436992 501190 437092
rect 501314 436992 501414 437092
rect 500418 436768 500518 436868
rect 500642 436768 500742 436868
rect 500866 436768 500966 436868
rect 501090 436768 501190 436868
rect 501314 436768 501414 436868
rect 500418 436544 500518 436644
rect 500642 436544 500742 436644
rect 500866 436544 500966 436644
rect 501090 436544 501190 436644
rect 501314 436544 501414 436644
rect 500418 436320 500518 436420
rect 500642 436320 500742 436420
rect 500866 436320 500966 436420
rect 501090 436320 501190 436420
rect 501314 436320 501414 436420
rect 500418 436096 500518 436196
rect 500642 436096 500742 436196
rect 500866 436096 500966 436196
rect 501090 436096 501190 436196
rect 501314 436096 501414 436196
rect 500418 435872 500518 435972
rect 500642 435872 500742 435972
rect 500866 435872 500966 435972
rect 501090 435872 501190 435972
rect 501314 435872 501414 435972
rect 500418 435648 500518 435748
rect 500642 435648 500742 435748
rect 500866 435648 500966 435748
rect 501090 435648 501190 435748
rect 501314 435648 501414 435748
rect 500418 435424 500518 435524
rect 500642 435424 500742 435524
rect 500866 435424 500966 435524
rect 501090 435424 501190 435524
rect 501314 435424 501414 435524
rect 500418 435200 500518 435300
rect 500642 435200 500742 435300
rect 500866 435200 500966 435300
rect 501090 435200 501190 435300
rect 501314 435200 501414 435300
rect 500418 434976 500518 435076
rect 500642 434976 500742 435076
rect 500866 434976 500966 435076
rect 501090 434976 501190 435076
rect 501314 434976 501414 435076
rect 512228 459336 513212 460204
rect 512228 457348 512422 459336
rect 512422 457348 512836 459336
rect 512836 457348 513212 459336
rect 512228 445636 513212 457348
rect 527618 460798 527718 460898
rect 527842 460798 527942 460898
rect 528066 460798 528166 460898
rect 528290 460798 528390 460898
rect 528514 460798 528614 460898
rect 527618 460574 527718 460674
rect 527842 460574 527942 460674
rect 528066 460574 528166 460674
rect 528290 460574 528390 460674
rect 528514 460574 528614 460674
rect 527618 460350 527718 460450
rect 527842 460350 527942 460450
rect 528066 460350 528166 460450
rect 528290 460350 528390 460450
rect 528514 460350 528614 460450
rect 527618 460126 527718 460226
rect 527842 460126 527942 460226
rect 528066 460126 528166 460226
rect 528290 460126 528390 460226
rect 528514 460126 528614 460226
rect 527618 459902 527718 460002
rect 527842 459902 527942 460002
rect 528066 459902 528166 460002
rect 528290 459902 528390 460002
rect 528514 459902 528614 460002
rect 527618 459678 527718 459778
rect 527842 459678 527942 459778
rect 528066 459678 528166 459778
rect 528290 459678 528390 459778
rect 528514 459678 528614 459778
rect 527618 459454 527718 459554
rect 527842 459454 527942 459554
rect 528066 459454 528166 459554
rect 528290 459454 528390 459554
rect 528514 459454 528614 459554
rect 527618 459230 527718 459330
rect 527842 459230 527942 459330
rect 528066 459230 528166 459330
rect 528290 459230 528390 459330
rect 528514 459230 528614 459330
rect 527618 459006 527718 459106
rect 527842 459006 527942 459106
rect 528066 459006 528166 459106
rect 528290 459006 528390 459106
rect 528514 459006 528614 459106
rect 527618 458782 527718 458882
rect 527842 458782 527942 458882
rect 528066 458782 528166 458882
rect 528290 458782 528390 458882
rect 528514 458782 528614 458882
rect 527618 458558 527718 458658
rect 527842 458558 527942 458658
rect 528066 458558 528166 458658
rect 528290 458558 528390 458658
rect 528514 458558 528614 458658
rect 527618 458334 527718 458434
rect 527842 458334 527942 458434
rect 528066 458334 528166 458434
rect 528290 458334 528390 458434
rect 528514 458334 528614 458434
rect 527618 458110 527718 458210
rect 527842 458110 527942 458210
rect 528066 458110 528166 458210
rect 528290 458110 528390 458210
rect 528514 458110 528614 458210
rect 527618 457886 527718 457986
rect 527842 457886 527942 457986
rect 528066 457886 528166 457986
rect 528290 457886 528390 457986
rect 528514 457886 528614 457986
rect 527618 457662 527718 457762
rect 527842 457662 527942 457762
rect 528066 457662 528166 457762
rect 528290 457662 528390 457762
rect 528514 457662 528614 457762
rect 527618 457438 527718 457538
rect 527842 457438 527942 457538
rect 528066 457438 528166 457538
rect 528290 457438 528390 457538
rect 528514 457438 528614 457538
rect 527618 457214 527718 457314
rect 527842 457214 527942 457314
rect 528066 457214 528166 457314
rect 528290 457214 528390 457314
rect 528514 457214 528614 457314
rect 562480 455360 562560 455440
rect 562640 455360 562720 455440
rect 562800 455360 562880 455440
rect 562960 455360 563040 455440
rect 563120 455360 563200 455440
rect 563280 455360 563360 455440
rect 563440 455360 563520 455440
rect 563600 455360 563680 455440
rect 563760 455360 563840 455440
rect 563920 455360 564000 455440
rect 564080 455360 564160 455440
rect 564240 455360 564320 455440
rect 564400 455360 564480 455440
rect 564560 455360 564640 455440
rect 564720 455360 564800 455440
rect 564880 455360 564960 455440
rect 565040 455360 565120 455440
rect 565200 455360 565280 455440
rect 565360 455360 565440 455440
rect 565520 455360 565600 455440
rect 565680 455360 565760 455440
rect 565840 455360 565920 455440
rect 566000 455360 566080 455440
rect 566160 455360 566240 455440
rect 566320 455360 566400 455440
rect 566480 455360 566560 455440
rect 566640 455360 566720 455440
rect 566800 455360 566880 455440
rect 566960 455360 567040 455440
rect 567120 455360 567200 455440
rect 567280 455360 567360 455440
rect 562480 455200 562560 455280
rect 562640 455200 562720 455280
rect 562800 455200 562880 455280
rect 562960 455200 563040 455280
rect 563120 455200 563200 455280
rect 563280 455200 563360 455280
rect 563440 455200 563520 455280
rect 563600 455200 563680 455280
rect 563760 455200 563840 455280
rect 563920 455200 564000 455280
rect 564080 455200 564160 455280
rect 564240 455200 564320 455280
rect 564400 455200 564480 455280
rect 564560 455200 564640 455280
rect 564720 455200 564800 455280
rect 564880 455200 564960 455280
rect 565040 455200 565120 455280
rect 565200 455200 565280 455280
rect 565360 455200 565440 455280
rect 565520 455200 565600 455280
rect 565680 455200 565760 455280
rect 565840 455200 565920 455280
rect 566000 455200 566080 455280
rect 566160 455200 566240 455280
rect 566320 455200 566400 455280
rect 566480 455200 566560 455280
rect 566640 455200 566720 455280
rect 566800 455200 566880 455280
rect 566960 455200 567040 455280
rect 567120 455200 567200 455280
rect 567280 455200 567360 455280
rect 572640 455360 572720 455440
rect 572800 455360 572880 455440
rect 572960 455360 573040 455440
rect 573120 455360 573200 455440
rect 573280 455360 573360 455440
rect 573440 455360 573520 455440
rect 573600 455360 573680 455440
rect 573760 455360 573840 455440
rect 573920 455360 574000 455440
rect 574080 455360 574160 455440
rect 574240 455360 574320 455440
rect 574400 455360 574480 455440
rect 574560 455360 574640 455440
rect 574720 455360 574800 455440
rect 574880 455360 574960 455440
rect 575040 455360 575120 455440
rect 575200 455360 575280 455440
rect 575360 455360 575440 455440
rect 575520 455360 575600 455440
rect 575680 455360 575760 455440
rect 575840 455360 575920 455440
rect 576000 455360 576080 455440
rect 576160 455360 576240 455440
rect 576320 455360 576400 455440
rect 576480 455360 576560 455440
rect 576640 455360 576720 455440
rect 576800 455360 576880 455440
rect 576960 455360 577040 455440
rect 577120 455360 577200 455440
rect 577280 455360 577360 455440
rect 577440 455360 577520 455440
rect 572640 455200 572720 455280
rect 572800 455200 572880 455280
rect 572960 455200 573040 455280
rect 573120 455200 573200 455280
rect 573280 455200 573360 455280
rect 573440 455200 573520 455280
rect 573600 455200 573680 455280
rect 573760 455200 573840 455280
rect 573920 455200 574000 455280
rect 574080 455200 574160 455280
rect 574240 455200 574320 455280
rect 574400 455200 574480 455280
rect 574560 455200 574640 455280
rect 574720 455200 574800 455280
rect 574880 455200 574960 455280
rect 575040 455200 575120 455280
rect 575200 455200 575280 455280
rect 575360 455200 575440 455280
rect 575520 455200 575600 455280
rect 575680 455200 575760 455280
rect 575840 455200 575920 455280
rect 576000 455200 576080 455280
rect 576160 455200 576240 455280
rect 576320 455200 576400 455280
rect 576480 455200 576560 455280
rect 576640 455200 576720 455280
rect 576800 455200 576880 455280
rect 576960 455200 577040 455280
rect 577120 455200 577200 455280
rect 577280 455200 577360 455280
rect 577440 455200 577520 455280
rect 562222 453859 562282 453919
rect 562342 453859 562402 453919
rect 562462 453859 562522 453919
rect 562582 453859 562642 453919
rect 562702 453859 562762 453919
rect 562822 453859 562882 453919
rect 562942 453859 563002 453919
rect 563062 453859 563122 453919
rect 563182 453859 563242 453919
rect 563302 453859 563362 453919
rect 563422 453859 563482 453919
rect 563542 453859 563602 453919
rect 563662 453859 563722 453919
rect 563782 453859 563842 453919
rect 563902 453859 563962 453919
rect 564022 453859 564082 453919
rect 564142 453859 564202 453919
rect 564262 453859 564322 453919
rect 564382 453859 564442 453919
rect 564502 453859 564562 453919
rect 564622 453859 564682 453919
rect 564742 453859 564802 453919
rect 564862 453859 564922 453919
rect 564982 453859 565042 453919
rect 565102 453859 565162 453919
rect 565222 453859 565282 453919
rect 565342 453859 565402 453919
rect 565462 453859 565522 453919
rect 565582 453859 565642 453919
rect 565702 453859 565762 453919
rect 565822 453859 565882 453919
rect 565942 453859 566002 453919
rect 566062 453859 566122 453919
rect 566182 453859 566242 453919
rect 566302 453859 566362 453919
rect 566422 453859 566482 453919
rect 566542 453859 566602 453919
rect 566662 453859 566722 453919
rect 566782 453859 566842 453919
rect 566902 453859 566962 453919
rect 567022 453859 567082 453919
rect 567142 453859 567202 453919
rect 567262 453859 567322 453919
rect 567382 453859 567442 453919
rect 567502 453859 567562 453919
rect 513720 453556 513920 453756
rect 514154 453556 514354 453756
rect 514588 453556 514788 453756
rect 562222 453739 562282 453799
rect 562342 453739 562402 453799
rect 562462 453739 562522 453799
rect 562582 453739 562642 453799
rect 562702 453739 562762 453799
rect 562822 453739 562882 453799
rect 562942 453739 563002 453799
rect 563062 453739 563122 453799
rect 563182 453739 563242 453799
rect 563302 453739 563362 453799
rect 563422 453739 563482 453799
rect 563542 453739 563602 453799
rect 563662 453739 563722 453799
rect 563782 453739 563842 453799
rect 563902 453739 563962 453799
rect 564022 453739 564082 453799
rect 564142 453739 564202 453799
rect 564262 453739 564322 453799
rect 564382 453739 564442 453799
rect 564502 453739 564562 453799
rect 564622 453739 564682 453799
rect 564742 453739 564802 453799
rect 564862 453739 564922 453799
rect 564982 453739 565042 453799
rect 565102 453739 565162 453799
rect 565222 453739 565282 453799
rect 565342 453739 565402 453799
rect 565462 453739 565522 453799
rect 565582 453739 565642 453799
rect 565702 453739 565762 453799
rect 565822 453739 565882 453799
rect 565942 453739 566002 453799
rect 566062 453739 566122 453799
rect 566182 453739 566242 453799
rect 566302 453739 566362 453799
rect 566422 453739 566482 453799
rect 566542 453739 566602 453799
rect 566662 453739 566722 453799
rect 566782 453739 566842 453799
rect 566902 453739 566962 453799
rect 567022 453739 567082 453799
rect 567142 453739 567202 453799
rect 567262 453739 567322 453799
rect 567382 453739 567442 453799
rect 567502 453739 567562 453799
rect 572332 453874 572392 453934
rect 572452 453874 572512 453934
rect 572572 453874 572632 453934
rect 572692 453874 572752 453934
rect 572812 453874 572872 453934
rect 572932 453874 572992 453934
rect 573052 453874 573112 453934
rect 573172 453874 573232 453934
rect 573292 453874 573352 453934
rect 573412 453874 573472 453934
rect 573532 453874 573592 453934
rect 573652 453874 573712 453934
rect 573772 453874 573832 453934
rect 573892 453874 573952 453934
rect 574012 453874 574072 453934
rect 574132 453874 574192 453934
rect 574252 453874 574312 453934
rect 574372 453874 574432 453934
rect 574492 453874 574552 453934
rect 574612 453874 574672 453934
rect 574732 453874 574792 453934
rect 574852 453874 574912 453934
rect 574972 453874 575032 453934
rect 575092 453874 575152 453934
rect 575212 453874 575272 453934
rect 575332 453874 575392 453934
rect 575452 453874 575512 453934
rect 575572 453874 575632 453934
rect 575692 453874 575752 453934
rect 575812 453874 575872 453934
rect 575932 453874 575992 453934
rect 576052 453874 576112 453934
rect 576172 453874 576232 453934
rect 576292 453874 576352 453934
rect 576412 453874 576472 453934
rect 576532 453874 576592 453934
rect 576652 453874 576712 453934
rect 576772 453874 576832 453934
rect 576892 453874 576952 453934
rect 577012 453874 577072 453934
rect 577132 453874 577192 453934
rect 577252 453874 577312 453934
rect 577372 453874 577432 453934
rect 577492 453874 577552 453934
rect 577612 453874 577672 453934
rect 572332 453754 572392 453814
rect 572452 453754 572512 453814
rect 572572 453754 572632 453814
rect 572692 453754 572752 453814
rect 572812 453754 572872 453814
rect 572932 453754 572992 453814
rect 573052 453754 573112 453814
rect 573172 453754 573232 453814
rect 573292 453754 573352 453814
rect 573412 453754 573472 453814
rect 573532 453754 573592 453814
rect 573652 453754 573712 453814
rect 573772 453754 573832 453814
rect 573892 453754 573952 453814
rect 574012 453754 574072 453814
rect 574132 453754 574192 453814
rect 574252 453754 574312 453814
rect 574372 453754 574432 453814
rect 574492 453754 574552 453814
rect 574612 453754 574672 453814
rect 574732 453754 574792 453814
rect 574852 453754 574912 453814
rect 574972 453754 575032 453814
rect 575092 453754 575152 453814
rect 575212 453754 575272 453814
rect 575332 453754 575392 453814
rect 575452 453754 575512 453814
rect 575572 453754 575632 453814
rect 575692 453754 575752 453814
rect 575812 453754 575872 453814
rect 575932 453754 575992 453814
rect 576052 453754 576112 453814
rect 576172 453754 576232 453814
rect 576292 453754 576352 453814
rect 576412 453754 576472 453814
rect 576532 453754 576592 453814
rect 576652 453754 576712 453814
rect 576772 453754 576832 453814
rect 576892 453754 576952 453814
rect 577012 453754 577072 453814
rect 577132 453754 577192 453814
rect 577252 453754 577312 453814
rect 577372 453754 577432 453814
rect 577492 453754 577552 453814
rect 577612 453754 577672 453814
rect 513720 453122 513920 453322
rect 514154 453122 514354 453322
rect 514588 453122 514788 453322
rect 513720 452688 513920 452888
rect 514154 452688 514354 452888
rect 514588 452688 514788 452888
rect 513720 452254 513920 452454
rect 514154 452254 514354 452454
rect 514588 452254 514788 452454
rect 513720 451820 513920 452020
rect 514154 451820 514354 452020
rect 514588 451820 514788 452020
rect 513720 451386 513920 451586
rect 514154 451386 514354 451586
rect 514588 451386 514788 451586
rect 513720 450952 513920 451152
rect 514154 450952 514354 451152
rect 514588 450952 514788 451152
rect 513720 450518 513920 450718
rect 514154 450518 514354 450718
rect 514588 450518 514788 450718
rect 513720 450084 513920 450284
rect 514154 450084 514354 450284
rect 514588 450084 514788 450284
rect 513720 449650 513920 449850
rect 514154 449650 514354 449850
rect 514588 449650 514788 449850
rect 513720 449216 513920 449416
rect 514154 449216 514354 449416
rect 514588 449216 514788 449416
rect 514588 448816 514788 449016
rect 514588 448416 514788 448616
rect 514588 448016 514788 448216
rect 514588 447616 514788 447816
rect 514588 447216 514788 447416
rect 514588 446816 514788 447016
rect 514588 446416 514788 446616
rect 514588 446016 514788 446216
rect 512228 443648 512422 445636
rect 512422 443648 512836 445636
rect 512836 443648 513212 445636
rect 514588 445616 514788 445816
rect 512228 440324 513212 443648
rect 514588 444016 514788 444216
rect 514588 443616 514788 443816
rect 514588 443216 514788 443416
rect 514588 442816 514788 443016
rect 514588 442416 514788 442616
rect 514588 442016 514788 442216
rect 514588 441616 514788 441816
rect 514588 441216 514788 441416
rect 514588 440816 514788 441016
rect 512228 439882 512836 440324
rect 512836 439882 513212 440324
rect 527638 437440 527738 437540
rect 527862 437440 527962 437540
rect 528086 437440 528186 437540
rect 528310 437440 528410 437540
rect 528534 437440 528634 437540
rect 527638 437216 527738 437316
rect 527862 437216 527962 437316
rect 528086 437216 528186 437316
rect 528310 437216 528410 437316
rect 528534 437216 528634 437316
rect 527638 436992 527738 437092
rect 527862 436992 527962 437092
rect 528086 436992 528186 437092
rect 528310 436992 528410 437092
rect 528534 436992 528634 437092
rect 527638 436768 527738 436868
rect 527862 436768 527962 436868
rect 528086 436768 528186 436868
rect 528310 436768 528410 436868
rect 528534 436768 528634 436868
rect 527638 436544 527738 436644
rect 527862 436544 527962 436644
rect 528086 436544 528186 436644
rect 528310 436544 528410 436644
rect 528534 436544 528634 436644
rect 527638 436320 527738 436420
rect 527862 436320 527962 436420
rect 528086 436320 528186 436420
rect 528310 436320 528410 436420
rect 528534 436320 528634 436420
rect 527638 436096 527738 436196
rect 527862 436096 527962 436196
rect 528086 436096 528186 436196
rect 528310 436096 528410 436196
rect 528534 436096 528634 436196
rect 527638 435872 527738 435972
rect 527862 435872 527962 435972
rect 528086 435872 528186 435972
rect 528310 435872 528410 435972
rect 528534 435872 528634 435972
rect 527638 435648 527738 435748
rect 527862 435648 527962 435748
rect 528086 435648 528186 435748
rect 528310 435648 528410 435748
rect 528534 435648 528634 435748
rect 527638 435424 527738 435524
rect 527862 435424 527962 435524
rect 528086 435424 528186 435524
rect 528310 435424 528410 435524
rect 528534 435424 528634 435524
rect 527638 435200 527738 435300
rect 527862 435200 527962 435300
rect 528086 435200 528186 435300
rect 528310 435200 528410 435300
rect 528534 435200 528634 435300
rect 527638 434976 527738 435076
rect 527862 434976 527962 435076
rect 528086 434976 528186 435076
rect 528310 434976 528410 435076
rect 528534 434976 528634 435076
rect 500418 434752 500518 434852
rect 500642 434752 500742 434852
rect 500866 434752 500966 434852
rect 501090 434752 501190 434852
rect 501314 434752 501414 434852
rect 500418 434528 500518 434628
rect 500642 434528 500742 434628
rect 500866 434528 500966 434628
rect 501090 434528 501190 434628
rect 501314 434528 501414 434628
rect 500418 434304 500518 434404
rect 500642 434304 500742 434404
rect 500866 434304 500966 434404
rect 501090 434304 501190 434404
rect 501314 434304 501414 434404
rect 500418 434080 500518 434180
rect 500642 434080 500742 434180
rect 500866 434080 500966 434180
rect 501090 434080 501190 434180
rect 501314 434080 501414 434180
rect 500418 433856 500518 433956
rect 500642 433856 500742 433956
rect 500866 433856 500966 433956
rect 501090 433856 501190 433956
rect 501314 433856 501414 433956
rect 500418 433632 500518 433732
rect 500642 433632 500742 433732
rect 500866 433632 500966 433732
rect 501090 433632 501190 433732
rect 501314 433632 501414 433732
rect 500418 433408 500518 433508
rect 500642 433408 500742 433508
rect 500866 433408 500966 433508
rect 501090 433408 501190 433508
rect 501314 433408 501414 433508
rect 500418 433184 500518 433284
rect 500642 433184 500742 433284
rect 500866 433184 500966 433284
rect 501090 433184 501190 433284
rect 501314 433184 501414 433284
rect 500418 432960 500518 433060
rect 500642 432960 500742 433060
rect 500866 432960 500966 433060
rect 501090 432960 501190 433060
rect 501314 432960 501414 433060
rect 500418 432736 500518 432836
rect 500642 432736 500742 432836
rect 500866 432736 500966 432836
rect 501090 432736 501190 432836
rect 501314 432736 501414 432836
rect 500418 432512 500518 432612
rect 500642 432512 500742 432612
rect 500866 432512 500966 432612
rect 501090 432512 501190 432612
rect 501314 432512 501414 432612
rect 500418 432288 500518 432388
rect 500642 432288 500742 432388
rect 500866 432288 500966 432388
rect 501090 432288 501190 432388
rect 501314 432288 501414 432388
rect 500418 432064 500518 432164
rect 500642 432064 500742 432164
rect 500866 432064 500966 432164
rect 501090 432064 501190 432164
rect 501314 432064 501414 432164
rect 500418 431840 500518 431940
rect 500642 431840 500742 431940
rect 500866 431840 500966 431940
rect 501090 431840 501190 431940
rect 501314 431840 501414 431940
rect 500418 431616 500518 431716
rect 500642 431616 500742 431716
rect 500866 431616 500966 431716
rect 501090 431616 501190 431716
rect 501314 431616 501414 431716
rect 500418 431392 500518 431492
rect 500642 431392 500742 431492
rect 500866 431392 500966 431492
rect 501090 431392 501190 431492
rect 501314 431392 501414 431492
rect 500418 431168 500518 431268
rect 500642 431168 500742 431268
rect 500866 431168 500966 431268
rect 501090 431168 501190 431268
rect 501314 431168 501414 431268
rect 527638 434752 527738 434852
rect 527862 434752 527962 434852
rect 528086 434752 528186 434852
rect 528310 434752 528410 434852
rect 528534 434752 528634 434852
rect 527638 434528 527738 434628
rect 527862 434528 527962 434628
rect 528086 434528 528186 434628
rect 528310 434528 528410 434628
rect 528534 434528 528634 434628
rect 527638 434304 527738 434404
rect 527862 434304 527962 434404
rect 528086 434304 528186 434404
rect 528310 434304 528410 434404
rect 528534 434304 528634 434404
rect 527638 434080 527738 434180
rect 527862 434080 527962 434180
rect 528086 434080 528186 434180
rect 528310 434080 528410 434180
rect 528534 434080 528634 434180
rect 527638 433856 527738 433956
rect 527862 433856 527962 433956
rect 528086 433856 528186 433956
rect 528310 433856 528410 433956
rect 528534 433856 528634 433956
rect 527638 433632 527738 433732
rect 527862 433632 527962 433732
rect 528086 433632 528186 433732
rect 528310 433632 528410 433732
rect 528534 433632 528634 433732
rect 527638 433408 527738 433508
rect 527862 433408 527962 433508
rect 528086 433408 528186 433508
rect 528310 433408 528410 433508
rect 528534 433408 528634 433508
rect 527638 433184 527738 433284
rect 527862 433184 527962 433284
rect 528086 433184 528186 433284
rect 528310 433184 528410 433284
rect 528534 433184 528634 433284
rect 527638 432960 527738 433060
rect 527862 432960 527962 433060
rect 528086 432960 528186 433060
rect 528310 432960 528410 433060
rect 528534 432960 528634 433060
rect 527638 432736 527738 432836
rect 527862 432736 527962 432836
rect 528086 432736 528186 432836
rect 528310 432736 528410 432836
rect 528534 432736 528634 432836
rect 527638 432512 527738 432612
rect 527862 432512 527962 432612
rect 528086 432512 528186 432612
rect 528310 432512 528410 432612
rect 528534 432512 528634 432612
rect 527638 432288 527738 432388
rect 527862 432288 527962 432388
rect 528086 432288 528186 432388
rect 528310 432288 528410 432388
rect 528534 432288 528634 432388
rect 527638 432064 527738 432164
rect 527862 432064 527962 432164
rect 528086 432064 528186 432164
rect 528310 432064 528410 432164
rect 528534 432064 528634 432164
rect 527638 431840 527738 431940
rect 527862 431840 527962 431940
rect 528086 431840 528186 431940
rect 528310 431840 528410 431940
rect 528534 431840 528634 431940
rect 527638 431616 527738 431716
rect 527862 431616 527962 431716
rect 528086 431616 528186 431716
rect 528310 431616 528410 431716
rect 528534 431616 528634 431716
rect 527638 431392 527738 431492
rect 527862 431392 527962 431492
rect 528086 431392 528186 431492
rect 528310 431392 528410 431492
rect 528534 431392 528634 431492
rect 527638 431168 527738 431268
rect 527862 431168 527962 431268
rect 528086 431168 528186 431268
rect 528310 431168 528410 431268
rect 528534 431168 528634 431268
rect 500418 430944 500518 431044
rect 500642 430944 500742 431044
rect 500866 430944 500966 431044
rect 501090 430944 501190 431044
rect 501314 430944 501414 431044
rect 503920 430926 504020 431026
rect 504144 430926 504244 431026
rect 504368 430926 504468 431026
rect 504592 430926 504692 431026
rect 504816 430926 504916 431026
rect 505040 430926 505140 431026
rect 505264 430926 505364 431026
rect 505488 430926 505588 431026
rect 505712 430926 505812 431026
rect 505936 430926 506036 431026
rect 506160 430926 506260 431026
rect 506384 430926 506484 431026
rect 506608 430926 506708 431026
rect 506832 430926 506932 431026
rect 507056 430926 507156 431026
rect 507280 430926 507380 431026
rect 507504 430926 507604 431026
rect 507728 430926 507828 431026
rect 507952 430926 508052 431026
rect 508176 430926 508276 431026
rect 508400 430926 508500 431026
rect 508624 430926 508724 431026
rect 508848 430926 508948 431026
rect 509072 430926 509172 431026
rect 509296 430926 509396 431026
rect 509520 430926 509620 431026
rect 509744 430926 509844 431026
rect 509968 430926 510068 431026
rect 510192 430926 510292 431026
rect 510416 430926 510516 431026
rect 503920 430702 504020 430802
rect 504144 430702 504244 430802
rect 504368 430702 504468 430802
rect 504592 430702 504692 430802
rect 504816 430702 504916 430802
rect 505040 430702 505140 430802
rect 505264 430702 505364 430802
rect 505488 430702 505588 430802
rect 505712 430702 505812 430802
rect 505936 430702 506036 430802
rect 506160 430702 506260 430802
rect 506384 430702 506484 430802
rect 506608 430702 506708 430802
rect 506832 430702 506932 430802
rect 507056 430702 507156 430802
rect 507280 430702 507380 430802
rect 507504 430702 507604 430802
rect 507728 430702 507828 430802
rect 507952 430702 508052 430802
rect 508176 430702 508276 430802
rect 508400 430702 508500 430802
rect 508624 430702 508724 430802
rect 508848 430702 508948 430802
rect 509072 430702 509172 430802
rect 509296 430702 509396 430802
rect 509520 430702 509620 430802
rect 509744 430702 509844 430802
rect 509968 430702 510068 430802
rect 510192 430702 510292 430802
rect 510416 430702 510516 430802
rect 503920 430478 504020 430578
rect 504144 430478 504244 430578
rect 504368 430478 504468 430578
rect 504592 430478 504692 430578
rect 504816 430478 504916 430578
rect 505040 430478 505140 430578
rect 505264 430478 505364 430578
rect 505488 430478 505588 430578
rect 505712 430478 505812 430578
rect 505936 430478 506036 430578
rect 506160 430478 506260 430578
rect 506384 430478 506484 430578
rect 506608 430478 506708 430578
rect 506832 430478 506932 430578
rect 507056 430478 507156 430578
rect 507280 430478 507380 430578
rect 507504 430478 507604 430578
rect 507728 430478 507828 430578
rect 507952 430478 508052 430578
rect 508176 430478 508276 430578
rect 508400 430478 508500 430578
rect 508624 430478 508724 430578
rect 508848 430478 508948 430578
rect 509072 430478 509172 430578
rect 509296 430478 509396 430578
rect 509520 430478 509620 430578
rect 509744 430478 509844 430578
rect 509968 430478 510068 430578
rect 510192 430478 510292 430578
rect 510416 430478 510516 430578
rect 503920 430254 504020 430354
rect 504144 430254 504244 430354
rect 504368 430254 504468 430354
rect 504592 430254 504692 430354
rect 504816 430254 504916 430354
rect 505040 430254 505140 430354
rect 505264 430254 505364 430354
rect 505488 430254 505588 430354
rect 505712 430254 505812 430354
rect 505936 430254 506036 430354
rect 506160 430254 506260 430354
rect 506384 430254 506484 430354
rect 506608 430254 506708 430354
rect 506832 430254 506932 430354
rect 507056 430254 507156 430354
rect 507280 430254 507380 430354
rect 507504 430254 507604 430354
rect 507728 430254 507828 430354
rect 507952 430254 508052 430354
rect 508176 430254 508276 430354
rect 508400 430254 508500 430354
rect 508624 430254 508724 430354
rect 508848 430254 508948 430354
rect 509072 430254 509172 430354
rect 509296 430254 509396 430354
rect 509520 430254 509620 430354
rect 509744 430254 509844 430354
rect 509968 430254 510068 430354
rect 510192 430254 510292 430354
rect 510416 430254 510516 430354
rect 503920 430030 504020 430130
rect 504144 430030 504244 430130
rect 504368 430030 504468 430130
rect 504592 430030 504692 430130
rect 504816 430030 504916 430130
rect 505040 430030 505140 430130
rect 505264 430030 505364 430130
rect 505488 430030 505588 430130
rect 505712 430030 505812 430130
rect 505936 430030 506036 430130
rect 506160 430030 506260 430130
rect 506384 430030 506484 430130
rect 506608 430030 506708 430130
rect 506832 430030 506932 430130
rect 507056 430030 507156 430130
rect 507280 430030 507380 430130
rect 507504 430030 507604 430130
rect 507728 430030 507828 430130
rect 507952 430030 508052 430130
rect 508176 430030 508276 430130
rect 508400 430030 508500 430130
rect 508624 430030 508724 430130
rect 508848 430030 508948 430130
rect 509072 430030 509172 430130
rect 509296 430030 509396 430130
rect 509520 430030 509620 430130
rect 509744 430030 509844 430130
rect 509968 430030 510068 430130
rect 510192 430030 510292 430130
rect 510416 430030 510516 430130
rect 517320 430926 517420 431026
rect 517544 430926 517644 431026
rect 517768 430926 517868 431026
rect 517992 430926 518092 431026
rect 518216 430926 518316 431026
rect 518440 430926 518540 431026
rect 518664 430926 518764 431026
rect 518888 430926 518988 431026
rect 519112 430926 519212 431026
rect 519336 430926 519436 431026
rect 519560 430926 519660 431026
rect 519784 430926 519884 431026
rect 520008 430926 520108 431026
rect 520232 430926 520332 431026
rect 520456 430926 520556 431026
rect 520680 430926 520780 431026
rect 520904 430926 521004 431026
rect 521128 430926 521228 431026
rect 521352 430926 521452 431026
rect 521576 430926 521676 431026
rect 521800 430926 521900 431026
rect 522024 430926 522124 431026
rect 522248 430926 522348 431026
rect 522472 430926 522572 431026
rect 522696 430926 522796 431026
rect 522920 430926 523020 431026
rect 523144 430926 523244 431026
rect 523368 430926 523468 431026
rect 523592 430926 523692 431026
rect 523816 430926 523916 431026
rect 527638 430944 527738 431044
rect 527862 430944 527962 431044
rect 528086 430944 528186 431044
rect 528310 430944 528410 431044
rect 528534 430944 528634 431044
rect 517320 430702 517420 430802
rect 517544 430702 517644 430802
rect 517768 430702 517868 430802
rect 517992 430702 518092 430802
rect 518216 430702 518316 430802
rect 518440 430702 518540 430802
rect 518664 430702 518764 430802
rect 518888 430702 518988 430802
rect 519112 430702 519212 430802
rect 519336 430702 519436 430802
rect 519560 430702 519660 430802
rect 519784 430702 519884 430802
rect 520008 430702 520108 430802
rect 520232 430702 520332 430802
rect 520456 430702 520556 430802
rect 520680 430702 520780 430802
rect 520904 430702 521004 430802
rect 521128 430702 521228 430802
rect 521352 430702 521452 430802
rect 521576 430702 521676 430802
rect 521800 430702 521900 430802
rect 522024 430702 522124 430802
rect 522248 430702 522348 430802
rect 522472 430702 522572 430802
rect 522696 430702 522796 430802
rect 522920 430702 523020 430802
rect 523144 430702 523244 430802
rect 523368 430702 523468 430802
rect 523592 430702 523692 430802
rect 523816 430702 523916 430802
rect 517320 430478 517420 430578
rect 517544 430478 517644 430578
rect 517768 430478 517868 430578
rect 517992 430478 518092 430578
rect 518216 430478 518316 430578
rect 518440 430478 518540 430578
rect 518664 430478 518764 430578
rect 518888 430478 518988 430578
rect 519112 430478 519212 430578
rect 519336 430478 519436 430578
rect 519560 430478 519660 430578
rect 519784 430478 519884 430578
rect 520008 430478 520108 430578
rect 520232 430478 520332 430578
rect 520456 430478 520556 430578
rect 520680 430478 520780 430578
rect 520904 430478 521004 430578
rect 521128 430478 521228 430578
rect 521352 430478 521452 430578
rect 521576 430478 521676 430578
rect 521800 430478 521900 430578
rect 522024 430478 522124 430578
rect 522248 430478 522348 430578
rect 522472 430478 522572 430578
rect 522696 430478 522796 430578
rect 522920 430478 523020 430578
rect 523144 430478 523244 430578
rect 523368 430478 523468 430578
rect 523592 430478 523692 430578
rect 523816 430478 523916 430578
rect 517320 430254 517420 430354
rect 517544 430254 517644 430354
rect 517768 430254 517868 430354
rect 517992 430254 518092 430354
rect 518216 430254 518316 430354
rect 518440 430254 518540 430354
rect 518664 430254 518764 430354
rect 518888 430254 518988 430354
rect 519112 430254 519212 430354
rect 519336 430254 519436 430354
rect 519560 430254 519660 430354
rect 519784 430254 519884 430354
rect 520008 430254 520108 430354
rect 520232 430254 520332 430354
rect 520456 430254 520556 430354
rect 520680 430254 520780 430354
rect 520904 430254 521004 430354
rect 521128 430254 521228 430354
rect 521352 430254 521452 430354
rect 521576 430254 521676 430354
rect 521800 430254 521900 430354
rect 522024 430254 522124 430354
rect 522248 430254 522348 430354
rect 522472 430254 522572 430354
rect 522696 430254 522796 430354
rect 522920 430254 523020 430354
rect 523144 430254 523244 430354
rect 523368 430254 523468 430354
rect 523592 430254 523692 430354
rect 523816 430254 523916 430354
rect 517320 430030 517420 430130
rect 517544 430030 517644 430130
rect 517768 430030 517868 430130
rect 517992 430030 518092 430130
rect 518216 430030 518316 430130
rect 518440 430030 518540 430130
rect 518664 430030 518764 430130
rect 518888 430030 518988 430130
rect 519112 430030 519212 430130
rect 519336 430030 519436 430130
rect 519560 430030 519660 430130
rect 519784 430030 519884 430130
rect 520008 430030 520108 430130
rect 520232 430030 520332 430130
rect 520456 430030 520556 430130
rect 520680 430030 520780 430130
rect 520904 430030 521004 430130
rect 521128 430030 521228 430130
rect 521352 430030 521452 430130
rect 521576 430030 521676 430130
rect 521800 430030 521900 430130
rect 522024 430030 522124 430130
rect 522248 430030 522348 430130
rect 522472 430030 522572 430130
rect 522696 430030 522796 430130
rect 522920 430030 523020 430130
rect 523144 430030 523244 430130
rect 523368 430030 523468 430130
rect 523592 430030 523692 430130
rect 523816 430030 523916 430130
<< metal3 >>
rect 16194 702300 21194 704800
rect 68194 702300 73194 704800
rect 120194 702300 125194 704800
rect 165594 702300 170594 704800
rect 170894 697200 173094 704800
rect 170894 692600 171000 697200
rect 173000 692600 173094 697200
rect 170894 692300 173094 692600
rect 173394 697200 175594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 173394 692600 173400 697200
rect 175400 692600 175594 697200
rect 173394 692300 175594 692600
rect 222594 697200 224794 704800
rect 222594 692600 222706 697200
rect 224706 692600 224794 697200
rect 222594 692300 224794 692600
rect 225094 697200 227294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 225094 692600 225106 697200
rect 227106 692600 227294 697200
rect 225094 692300 227294 692600
rect 324294 697200 326494 704800
rect 324294 692600 324412 697200
rect 326412 692600 326494 697200
rect 324294 692300 326494 692600
rect 326794 697200 328994 704800
rect 329294 702300 334294 704800
rect 413394 702300 418394 704800
rect 465394 702400 470394 704800
rect 326794 692600 326812 697200
rect 328812 692600 328994 697200
rect 326794 692300 328994 692600
rect 510594 697360 515394 704800
rect 510594 692560 510654 697360
rect 515334 692560 515394 697360
rect 510594 692500 515394 692560
rect 520594 697360 525394 704800
rect 566594 697380 571594 704800
rect 520594 692560 520654 697360
rect 525334 692560 525394 697360
rect 520594 692500 525394 692560
rect -800 680242 1700 685242
rect 577380 677984 584800 682984
rect -800 643842 1660 648642
rect 562480 644524 584800 644584
rect 562480 639844 562600 644524
rect 567400 639844 584800 644524
rect 562480 639784 584800 639844
rect -800 633842 1660 638642
rect 562540 634524 584800 634584
rect 562540 629844 562600 634524
rect 567400 629844 584800 634524
rect 562540 629784 584800 629844
rect 583520 589472 584800 589584
rect 583520 588290 584800 588402
rect 583520 587108 584800 587220
rect 583520 585926 584800 586038
rect 583520 584744 584800 584856
rect 583520 583562 584800 583674
rect -800 559442 1660 564242
rect -800 549442 1660 554242
rect 582340 550562 584800 555362
rect 582340 540562 584800 545362
rect 477192 522892 483800 523098
rect 562388 522892 567660 523006
rect 477060 522862 567660 522892
rect 477060 522626 477192 522862
rect 477428 522626 477664 522862
rect 477900 522626 478136 522862
rect 478372 522626 478608 522862
rect 478844 522626 479080 522862
rect 479316 522626 479552 522862
rect 479788 522626 480024 522862
rect 480260 522626 480496 522862
rect 480732 522626 480968 522862
rect 481204 522626 481440 522862
rect 481676 522626 481912 522862
rect 482148 522626 482384 522862
rect 482620 522626 482856 522862
rect 483092 522626 483328 522862
rect 483564 522740 567660 522862
rect 483564 522626 562624 522740
rect 477060 522504 562624 522626
rect 562860 522504 563096 522740
rect 563332 522504 563568 522740
rect 563804 522504 564040 522740
rect 564276 522504 564512 522740
rect 564748 522504 564984 522740
rect 565220 522504 565456 522740
rect 565692 522504 565928 522740
rect 566164 522504 566400 522740
rect 566636 522504 566872 522740
rect 567108 522504 567660 522740
rect 477060 522390 567660 522504
rect 477060 522154 477192 522390
rect 477428 522154 477664 522390
rect 477900 522154 478136 522390
rect 478372 522154 478608 522390
rect 478844 522154 479080 522390
rect 479316 522154 479552 522390
rect 479788 522154 480024 522390
rect 480260 522154 480496 522390
rect 480732 522154 480968 522390
rect 481204 522154 481440 522390
rect 481676 522154 481912 522390
rect 482148 522154 482384 522390
rect 482620 522154 482856 522390
rect 483092 522154 483328 522390
rect 483564 522268 567660 522390
rect 483564 522154 562624 522268
rect 477060 522032 562624 522154
rect 562860 522032 563096 522268
rect 563332 522032 563568 522268
rect 563804 522032 564040 522268
rect 564276 522032 564512 522268
rect 564748 522032 564984 522268
rect 565220 522032 565456 522268
rect 565692 522032 565928 522268
rect 566164 522032 566400 522268
rect 566636 522032 566872 522268
rect 567108 522032 567660 522268
rect 477060 521918 567660 522032
rect 477060 521682 477192 521918
rect 477428 521682 477664 521918
rect 477900 521682 478136 521918
rect 478372 521682 478608 521918
rect 478844 521682 479080 521918
rect 479316 521682 479552 521918
rect 479788 521682 480024 521918
rect 480260 521682 480496 521918
rect 480732 521682 480968 521918
rect 481204 521682 481440 521918
rect 481676 521682 481912 521918
rect 482148 521682 482384 521918
rect 482620 521682 482856 521918
rect 483092 521682 483328 521918
rect 483564 521796 567660 521918
rect 483564 521682 562624 521796
rect 477060 521560 562624 521682
rect 562860 521560 563096 521796
rect 563332 521560 563568 521796
rect 563804 521560 564040 521796
rect 564276 521560 564512 521796
rect 564748 521560 564984 521796
rect 565220 521560 565456 521796
rect 565692 521560 565928 521796
rect 566164 521560 566400 521796
rect 566636 521560 566872 521796
rect 567108 521560 567660 521796
rect 477060 521446 567660 521560
rect 477060 521210 477192 521446
rect 477428 521210 477664 521446
rect 477900 521210 478136 521446
rect 478372 521210 478608 521446
rect 478844 521210 479080 521446
rect 479316 521210 479552 521446
rect 479788 521210 480024 521446
rect 480260 521210 480496 521446
rect 480732 521210 480968 521446
rect 481204 521210 481440 521446
rect 481676 521210 481912 521446
rect 482148 521210 482384 521446
rect 482620 521210 482856 521446
rect 483092 521210 483328 521446
rect 483564 521324 567660 521446
rect 483564 521210 562624 521324
rect 477060 521088 562624 521210
rect 562860 521088 563096 521324
rect 563332 521088 563568 521324
rect 563804 521088 564040 521324
rect 564276 521088 564512 521324
rect 564748 521088 564984 521324
rect 565220 521088 565456 521324
rect 565692 521088 565928 521324
rect 566164 521088 566400 521324
rect 566636 521088 566872 521324
rect 567108 521088 567660 521324
rect 477060 520974 567660 521088
rect 477060 520738 477192 520974
rect 477428 520738 477664 520974
rect 477900 520738 478136 520974
rect 478372 520738 478608 520974
rect 478844 520738 479080 520974
rect 479316 520738 479552 520974
rect 479788 520738 480024 520974
rect 480260 520738 480496 520974
rect 480732 520738 480968 520974
rect 481204 520738 481440 520974
rect 481676 520738 481912 520974
rect 482148 520738 482384 520974
rect 482620 520738 482856 520974
rect 483092 520738 483328 520974
rect 483564 520852 567660 520974
rect 483564 520738 562624 520852
rect 477060 520616 562624 520738
rect 562860 520616 563096 520852
rect 563332 520616 563568 520852
rect 563804 520616 564040 520852
rect 564276 520616 564512 520852
rect 564748 520616 564984 520852
rect 565220 520616 565456 520852
rect 565692 520616 565928 520852
rect 566164 520616 566400 520852
rect 566636 520616 566872 520852
rect 567108 520616 567660 520852
rect 477060 520502 567660 520616
rect 477060 520266 477192 520502
rect 477428 520266 477664 520502
rect 477900 520266 478136 520502
rect 478372 520266 478608 520502
rect 478844 520266 479080 520502
rect 479316 520266 479552 520502
rect 479788 520266 480024 520502
rect 480260 520266 480496 520502
rect 480732 520266 480968 520502
rect 481204 520266 481440 520502
rect 481676 520266 481912 520502
rect 482148 520266 482384 520502
rect 482620 520266 482856 520502
rect 483092 520266 483328 520502
rect 483564 520380 567660 520502
rect 483564 520266 562624 520380
rect 477060 520144 562624 520266
rect 562860 520144 563096 520380
rect 563332 520144 563568 520380
rect 563804 520144 564040 520380
rect 564276 520144 564512 520380
rect 564748 520144 564984 520380
rect 565220 520144 565456 520380
rect 565692 520144 565928 520380
rect 566164 520144 566400 520380
rect 566636 520144 566872 520380
rect 567108 520144 567660 520380
rect 477060 520030 567660 520144
rect 477060 519794 477192 520030
rect 477428 519794 477664 520030
rect 477900 519794 478136 520030
rect 478372 519794 478608 520030
rect 478844 519794 479080 520030
rect 479316 519794 479552 520030
rect 479788 519794 480024 520030
rect 480260 519794 480496 520030
rect 480732 519794 480968 520030
rect 481204 519794 481440 520030
rect 481676 519794 481912 520030
rect 482148 519794 482384 520030
rect 482620 519794 482856 520030
rect 483092 519794 483328 520030
rect 483564 519908 567660 520030
rect 483564 519794 562624 519908
rect 477060 519672 562624 519794
rect 562860 519672 563096 519908
rect 563332 519672 563568 519908
rect 563804 519672 564040 519908
rect 564276 519672 564512 519908
rect 564748 519672 564984 519908
rect 565220 519672 565456 519908
rect 565692 519672 565928 519908
rect 566164 519672 566400 519908
rect 566636 519672 566872 519908
rect 567108 519672 567660 519908
rect 477060 519558 567660 519672
rect 477060 519322 477192 519558
rect 477428 519322 477664 519558
rect 477900 519322 478136 519558
rect 478372 519322 478608 519558
rect 478844 519322 479080 519558
rect 479316 519322 479552 519558
rect 479788 519322 480024 519558
rect 480260 519322 480496 519558
rect 480732 519322 480968 519558
rect 481204 519322 481440 519558
rect 481676 519322 481912 519558
rect 482148 519322 482384 519558
rect 482620 519322 482856 519558
rect 483092 519322 483328 519558
rect 483564 519436 567660 519558
rect 483564 519322 562624 519436
rect 477060 519200 562624 519322
rect 562860 519200 563096 519436
rect 563332 519200 563568 519436
rect 563804 519200 564040 519436
rect 564276 519200 564512 519436
rect 564748 519200 564984 519436
rect 565220 519200 565456 519436
rect 565692 519200 565928 519436
rect 566164 519200 566400 519436
rect 566636 519200 566872 519436
rect 567108 519200 567660 519436
rect 477060 519086 567660 519200
rect 477060 518850 477192 519086
rect 477428 518850 477664 519086
rect 477900 518850 478136 519086
rect 478372 518850 478608 519086
rect 478844 518850 479080 519086
rect 479316 518850 479552 519086
rect 479788 518850 480024 519086
rect 480260 518850 480496 519086
rect 480732 518850 480968 519086
rect 481204 518850 481440 519086
rect 481676 518850 481912 519086
rect 482148 518850 482384 519086
rect 482620 518850 482856 519086
rect 483092 518850 483328 519086
rect 483564 518964 567660 519086
rect 483564 518850 562624 518964
rect 477060 518728 562624 518850
rect 562860 518728 563096 518964
rect 563332 518728 563568 518964
rect 563804 518728 564040 518964
rect 564276 518728 564512 518964
rect 564748 518728 564984 518964
rect 565220 518728 565456 518964
rect 565692 518728 565928 518964
rect 566164 518728 566400 518964
rect 566636 518728 566872 518964
rect 567108 518728 567660 518964
rect 477060 518614 567660 518728
rect 477060 518378 477192 518614
rect 477428 518378 477664 518614
rect 477900 518378 478136 518614
rect 478372 518378 478608 518614
rect 478844 518378 479080 518614
rect 479316 518378 479552 518614
rect 479788 518378 480024 518614
rect 480260 518378 480496 518614
rect 480732 518378 480968 518614
rect 481204 518378 481440 518614
rect 481676 518378 481912 518614
rect 482148 518378 482384 518614
rect 482620 518378 482856 518614
rect 483092 518378 483328 518614
rect 483564 518492 567660 518614
rect 483564 518378 562624 518492
rect 477060 518256 562624 518378
rect 562860 518256 563096 518492
rect 563332 518256 563568 518492
rect 563804 518256 564040 518492
rect 564276 518256 564512 518492
rect 564748 518256 564984 518492
rect 565220 518256 565456 518492
rect 565692 518256 565928 518492
rect 566164 518256 566400 518492
rect 566636 518256 566872 518492
rect 567108 518256 567660 518492
rect 477060 518142 567660 518256
rect 477060 517906 477192 518142
rect 477428 517906 477664 518142
rect 477900 517906 478136 518142
rect 478372 517906 478608 518142
rect 478844 517906 479080 518142
rect 479316 517906 479552 518142
rect 479788 517906 480024 518142
rect 480260 517906 480496 518142
rect 480732 517906 480968 518142
rect 481204 517906 481440 518142
rect 481676 517906 481912 518142
rect 482148 517906 482384 518142
rect 482620 517906 482856 518142
rect 483092 517906 483328 518142
rect 483564 518020 567660 518142
rect 483564 517906 562624 518020
rect 477060 517784 562624 517906
rect 562860 517784 563096 518020
rect 563332 517784 563568 518020
rect 563804 517784 564040 518020
rect 564276 517784 564512 518020
rect 564748 517784 564984 518020
rect 565220 517784 565456 518020
rect 565692 517784 565928 518020
rect 566164 517784 566400 518020
rect 566636 517784 566872 518020
rect 567108 517784 567660 518020
rect 477060 517670 567660 517784
rect 477060 517434 477192 517670
rect 477428 517434 477664 517670
rect 477900 517434 478136 517670
rect 478372 517434 478608 517670
rect 478844 517434 479080 517670
rect 479316 517434 479552 517670
rect 479788 517434 480024 517670
rect 480260 517434 480496 517670
rect 480732 517434 480968 517670
rect 481204 517434 481440 517670
rect 481676 517434 481912 517670
rect 482148 517434 482384 517670
rect 482620 517434 482856 517670
rect 483092 517434 483328 517670
rect 483564 517548 567660 517670
rect 483564 517434 562624 517548
rect 477060 517312 562624 517434
rect 562860 517312 563096 517548
rect 563332 517312 563568 517548
rect 563804 517312 564040 517548
rect 564276 517312 564512 517548
rect 564748 517312 564984 517548
rect 565220 517312 565456 517548
rect 565692 517312 565928 517548
rect 566164 517312 566400 517548
rect 566636 517312 566872 517548
rect 567108 517312 567660 517548
rect 477060 517198 567660 517312
rect 477060 516962 477192 517198
rect 477428 516962 477664 517198
rect 477900 516962 478136 517198
rect 478372 516962 478608 517198
rect 478844 516962 479080 517198
rect 479316 516962 479552 517198
rect 479788 516962 480024 517198
rect 480260 516962 480496 517198
rect 480732 516962 480968 517198
rect 481204 516962 481440 517198
rect 481676 516962 481912 517198
rect 482148 516962 482384 517198
rect 482620 516962 482856 517198
rect 483092 516962 483328 517198
rect 483564 517076 567660 517198
rect 483564 516962 562624 517076
rect 477060 516840 562624 516962
rect 562860 516840 563096 517076
rect 563332 516840 563568 517076
rect 563804 516840 564040 517076
rect 564276 516840 564512 517076
rect 564748 516840 564984 517076
rect 565220 516840 565456 517076
rect 565692 516840 565928 517076
rect 566164 516840 566400 517076
rect 566636 516840 566872 517076
rect 567108 516840 567660 517076
rect 477060 516726 567660 516840
rect 477060 516490 477192 516726
rect 477428 516490 477664 516726
rect 477900 516490 478136 516726
rect 478372 516490 478608 516726
rect 478844 516490 479080 516726
rect 479316 516490 479552 516726
rect 479788 516490 480024 516726
rect 480260 516490 480496 516726
rect 480732 516490 480968 516726
rect 481204 516490 481440 516726
rect 481676 516490 481912 516726
rect 482148 516490 482384 516726
rect 482620 516490 482856 516726
rect 483092 516490 483328 516726
rect 483564 516604 567660 516726
rect 483564 516490 562624 516604
rect 477060 516368 562624 516490
rect 562860 516368 563096 516604
rect 563332 516368 563568 516604
rect 563804 516368 564040 516604
rect 564276 516368 564512 516604
rect 564748 516368 564984 516604
rect 565220 516368 565456 516604
rect 565692 516368 565928 516604
rect 566164 516368 566400 516604
rect 566636 516368 566872 516604
rect 567108 516368 567660 516604
rect 477060 516226 567660 516368
rect -800 511530 480 511642
rect -800 510348 480 510460
rect -800 509166 480 509278
rect -800 507984 480 508096
rect -800 506802 480 506914
rect -800 505620 480 505732
rect 583520 500050 584800 500162
rect 583520 498868 584800 498980
rect 583520 497686 584800 497798
rect 583520 496504 584800 496616
rect 562380 495742 567480 495822
rect 562380 495662 562480 495742
rect 562560 495662 562640 495742
rect 562720 495662 562800 495742
rect 562880 495662 562960 495742
rect 563040 495662 563120 495742
rect 563200 495662 563280 495742
rect 563360 495662 563440 495742
rect 563520 495662 563600 495742
rect 563680 495662 563760 495742
rect 563840 495662 563920 495742
rect 564000 495662 564080 495742
rect 564160 495662 564240 495742
rect 564320 495662 564400 495742
rect 564480 495662 564560 495742
rect 564640 495662 564720 495742
rect 564800 495662 564880 495742
rect 564960 495662 565040 495742
rect 565120 495662 565200 495742
rect 565280 495662 565360 495742
rect 565440 495662 565520 495742
rect 565600 495662 565680 495742
rect 565760 495662 565840 495742
rect 565920 495662 566000 495742
rect 566080 495662 566160 495742
rect 566240 495662 566320 495742
rect 566400 495662 566480 495742
rect 566560 495662 566640 495742
rect 566720 495662 566800 495742
rect 566880 495662 566960 495742
rect 567040 495662 567120 495742
rect 567200 495662 567280 495742
rect 567360 495662 567480 495742
rect 562380 495582 567480 495662
rect 562380 495502 562480 495582
rect 562560 495502 562640 495582
rect 562720 495502 562800 495582
rect 562880 495502 562960 495582
rect 563040 495502 563120 495582
rect 563200 495502 563280 495582
rect 563360 495502 563440 495582
rect 563520 495502 563600 495582
rect 563680 495502 563760 495582
rect 563840 495502 563920 495582
rect 564000 495502 564080 495582
rect 564160 495502 564240 495582
rect 564320 495502 564400 495582
rect 564480 495502 564560 495582
rect 564640 495502 564720 495582
rect 564800 495502 564880 495582
rect 564960 495502 565040 495582
rect 565120 495502 565200 495582
rect 565280 495502 565360 495582
rect 565440 495502 565520 495582
rect 565600 495502 565680 495582
rect 565760 495502 565840 495582
rect 565920 495502 566000 495582
rect 566080 495502 566160 495582
rect 566240 495502 566320 495582
rect 566400 495502 566480 495582
rect 566560 495502 566640 495582
rect 566720 495502 566800 495582
rect 566880 495502 566960 495582
rect 567040 495502 567120 495582
rect 567200 495502 567280 495582
rect 567360 495502 567480 495582
rect 562380 495462 567480 495502
rect 572540 495742 577640 495822
rect 572540 495662 572640 495742
rect 572720 495662 572800 495742
rect 572880 495662 572960 495742
rect 573040 495662 573120 495742
rect 573200 495662 573280 495742
rect 573360 495662 573440 495742
rect 573520 495662 573600 495742
rect 573680 495662 573760 495742
rect 573840 495662 573920 495742
rect 574000 495662 574080 495742
rect 574160 495662 574240 495742
rect 574320 495662 574400 495742
rect 574480 495662 574560 495742
rect 574640 495662 574720 495742
rect 574800 495662 574880 495742
rect 574960 495662 575040 495742
rect 575120 495662 575200 495742
rect 575280 495662 575360 495742
rect 575440 495662 575520 495742
rect 575600 495662 575680 495742
rect 575760 495662 575840 495742
rect 575920 495662 576000 495742
rect 576080 495662 576160 495742
rect 576240 495662 576320 495742
rect 576400 495662 576480 495742
rect 576560 495662 576640 495742
rect 576720 495662 576800 495742
rect 576880 495662 576960 495742
rect 577040 495662 577120 495742
rect 577200 495662 577280 495742
rect 577360 495662 577440 495742
rect 577520 495662 577640 495742
rect 572540 495582 577640 495662
rect 572540 495502 572640 495582
rect 572720 495502 572800 495582
rect 572880 495502 572960 495582
rect 573040 495502 573120 495582
rect 573200 495502 573280 495582
rect 573360 495502 573440 495582
rect 573520 495502 573600 495582
rect 573680 495502 573760 495582
rect 573840 495502 573920 495582
rect 574000 495502 574080 495582
rect 574160 495502 574240 495582
rect 574320 495502 574400 495582
rect 574480 495502 574560 495582
rect 574640 495502 574720 495582
rect 574800 495502 574880 495582
rect 574960 495502 575040 495582
rect 575120 495502 575200 495582
rect 575280 495502 575360 495582
rect 575440 495502 575520 495582
rect 575600 495502 575680 495582
rect 575760 495502 575840 495582
rect 575920 495502 576000 495582
rect 576080 495502 576160 495582
rect 576240 495502 576320 495582
rect 576400 495502 576480 495582
rect 576560 495502 576640 495582
rect 576720 495502 576800 495582
rect 576880 495502 576960 495582
rect 577040 495502 577120 495582
rect 577200 495502 577280 495582
rect 577360 495502 577440 495582
rect 577520 495502 577640 495582
rect 572540 495462 577640 495502
rect 583520 495322 584800 495434
rect 511400 494528 583800 494600
rect 511400 494464 511616 494528
rect 511680 494464 511744 494528
rect 511808 494464 511872 494528
rect 511936 494464 512000 494528
rect 512064 494464 583800 494528
rect 511400 494400 583800 494464
rect 511400 494336 511616 494400
rect 511680 494336 511744 494400
rect 511808 494336 511872 494400
rect 511936 494336 512000 494400
rect 512064 494336 583800 494400
rect 511400 494272 583800 494336
rect 511400 494208 511616 494272
rect 511680 494208 511744 494272
rect 511808 494208 511872 494272
rect 511936 494208 512000 494272
rect 512064 494252 583800 494272
rect 512064 494236 584800 494252
rect 512064 494221 572332 494236
rect 512064 494208 562222 494221
rect 511400 494161 562222 494208
rect 562282 494161 562342 494221
rect 562402 494161 562462 494221
rect 562522 494161 562582 494221
rect 562642 494161 562702 494221
rect 562762 494161 562822 494221
rect 562882 494161 562942 494221
rect 563002 494161 563062 494221
rect 563122 494161 563182 494221
rect 563242 494161 563302 494221
rect 563362 494161 563422 494221
rect 563482 494161 563542 494221
rect 563602 494161 563662 494221
rect 563722 494161 563782 494221
rect 563842 494161 563902 494221
rect 563962 494161 564022 494221
rect 564082 494161 564142 494221
rect 564202 494161 564262 494221
rect 564322 494161 564382 494221
rect 564442 494161 564502 494221
rect 564562 494161 564622 494221
rect 564682 494161 564742 494221
rect 564802 494161 564862 494221
rect 564922 494161 564982 494221
rect 565042 494161 565102 494221
rect 565162 494161 565222 494221
rect 565282 494161 565342 494221
rect 565402 494161 565462 494221
rect 565522 494161 565582 494221
rect 565642 494161 565702 494221
rect 565762 494161 565822 494221
rect 565882 494161 565942 494221
rect 566002 494161 566062 494221
rect 566122 494161 566182 494221
rect 566242 494161 566302 494221
rect 566362 494161 566422 494221
rect 566482 494161 566542 494221
rect 566602 494161 566662 494221
rect 566722 494161 566782 494221
rect 566842 494161 566902 494221
rect 566962 494161 567022 494221
rect 567082 494161 567142 494221
rect 567202 494161 567262 494221
rect 567322 494161 567382 494221
rect 567442 494161 567502 494221
rect 567562 494176 572332 494221
rect 572392 494176 572452 494236
rect 572512 494176 572572 494236
rect 572632 494176 572692 494236
rect 572752 494176 572812 494236
rect 572872 494176 572932 494236
rect 572992 494176 573052 494236
rect 573112 494176 573172 494236
rect 573232 494176 573292 494236
rect 573352 494176 573412 494236
rect 573472 494176 573532 494236
rect 573592 494176 573652 494236
rect 573712 494176 573772 494236
rect 573832 494176 573892 494236
rect 573952 494176 574012 494236
rect 574072 494176 574132 494236
rect 574192 494176 574252 494236
rect 574312 494176 574372 494236
rect 574432 494176 574492 494236
rect 574552 494176 574612 494236
rect 574672 494176 574732 494236
rect 574792 494176 574852 494236
rect 574912 494176 574972 494236
rect 575032 494176 575092 494236
rect 575152 494176 575212 494236
rect 575272 494176 575332 494236
rect 575392 494176 575452 494236
rect 575512 494176 575572 494236
rect 575632 494176 575692 494236
rect 575752 494176 575812 494236
rect 575872 494176 575932 494236
rect 575992 494176 576052 494236
rect 576112 494176 576172 494236
rect 576232 494176 576292 494236
rect 576352 494176 576412 494236
rect 576472 494176 576532 494236
rect 576592 494176 576652 494236
rect 576712 494176 576772 494236
rect 576832 494176 576892 494236
rect 576952 494176 577012 494236
rect 577072 494176 577132 494236
rect 577192 494176 577252 494236
rect 577312 494176 577372 494236
rect 577432 494176 577492 494236
rect 577552 494176 577612 494236
rect 577672 494176 584800 494236
rect 567562 494161 584800 494176
rect 511400 494144 584800 494161
rect 511400 494080 511616 494144
rect 511680 494080 511744 494144
rect 511808 494080 511872 494144
rect 511936 494080 512000 494144
rect 512064 494140 584800 494144
rect 512064 494116 583800 494140
rect 512064 494101 572332 494116
rect 512064 494080 562222 494101
rect 511400 494041 562222 494080
rect 562282 494041 562342 494101
rect 562402 494041 562462 494101
rect 562522 494041 562582 494101
rect 562642 494041 562702 494101
rect 562762 494041 562822 494101
rect 562882 494041 562942 494101
rect 563002 494041 563062 494101
rect 563122 494041 563182 494101
rect 563242 494041 563302 494101
rect 563362 494041 563422 494101
rect 563482 494041 563542 494101
rect 563602 494041 563662 494101
rect 563722 494041 563782 494101
rect 563842 494041 563902 494101
rect 563962 494041 564022 494101
rect 564082 494041 564142 494101
rect 564202 494041 564262 494101
rect 564322 494041 564382 494101
rect 564442 494041 564502 494101
rect 564562 494041 564622 494101
rect 564682 494041 564742 494101
rect 564802 494041 564862 494101
rect 564922 494041 564982 494101
rect 565042 494041 565102 494101
rect 565162 494041 565222 494101
rect 565282 494041 565342 494101
rect 565402 494041 565462 494101
rect 565522 494041 565582 494101
rect 565642 494041 565702 494101
rect 565762 494041 565822 494101
rect 565882 494041 565942 494101
rect 566002 494041 566062 494101
rect 566122 494041 566182 494101
rect 566242 494041 566302 494101
rect 566362 494041 566422 494101
rect 566482 494041 566542 494101
rect 566602 494041 566662 494101
rect 566722 494041 566782 494101
rect 566842 494041 566902 494101
rect 566962 494041 567022 494101
rect 567082 494041 567142 494101
rect 567202 494041 567262 494101
rect 567322 494041 567382 494101
rect 567442 494041 567502 494101
rect 567562 494056 572332 494101
rect 572392 494056 572452 494116
rect 572512 494056 572572 494116
rect 572632 494056 572692 494116
rect 572752 494056 572812 494116
rect 572872 494056 572932 494116
rect 572992 494056 573052 494116
rect 573112 494056 573172 494116
rect 573232 494056 573292 494116
rect 573352 494056 573412 494116
rect 573472 494056 573532 494116
rect 573592 494056 573652 494116
rect 573712 494056 573772 494116
rect 573832 494056 573892 494116
rect 573952 494056 574012 494116
rect 574072 494056 574132 494116
rect 574192 494056 574252 494116
rect 574312 494056 574372 494116
rect 574432 494056 574492 494116
rect 574552 494056 574612 494116
rect 574672 494056 574732 494116
rect 574792 494056 574852 494116
rect 574912 494056 574972 494116
rect 575032 494056 575092 494116
rect 575152 494056 575212 494116
rect 575272 494056 575332 494116
rect 575392 494056 575452 494116
rect 575512 494056 575572 494116
rect 575632 494056 575692 494116
rect 575752 494056 575812 494116
rect 575872 494056 575932 494116
rect 575992 494056 576052 494116
rect 576112 494056 576172 494116
rect 576232 494056 576292 494116
rect 576352 494056 576412 494116
rect 576472 494056 576532 494116
rect 576592 494056 576652 494116
rect 576712 494056 576772 494116
rect 576832 494056 576892 494116
rect 576952 494056 577012 494116
rect 577072 494056 577132 494116
rect 577192 494056 577252 494116
rect 577312 494056 577372 494116
rect 577432 494056 577492 494116
rect 577552 494056 577612 494116
rect 577672 494056 583800 494116
rect 567562 494041 583800 494056
rect 511400 494016 583800 494041
rect 511400 493952 511616 494016
rect 511680 493952 511744 494016
rect 511808 493952 511872 494016
rect 511936 493952 512000 494016
rect 512064 493952 583800 494016
rect 511400 493888 583800 493952
rect 511400 493824 511616 493888
rect 511680 493824 511744 493888
rect 511808 493824 511872 493888
rect 511936 493824 512000 493888
rect 512064 493824 583800 493888
rect 511400 493800 583800 493824
rect 572536 484236 577492 484272
rect 490440 483800 578504 484236
rect 490440 483564 572772 483800
rect 573008 483564 573244 483800
rect 573480 483564 573716 483800
rect 573952 483564 574188 483800
rect 574424 483564 574660 483800
rect 574896 483564 575132 483800
rect 575368 483564 575604 483800
rect 575840 483564 576076 483800
rect 576312 483564 576548 483800
rect 576784 483564 577020 483800
rect 577256 483564 578504 483800
rect 490440 483328 578504 483564
rect 490440 483236 572772 483328
rect 490440 478452 490940 483236
rect 496684 478452 503960 483236
rect 509704 478452 517360 483236
rect 523104 478452 530760 483236
rect 536504 483092 572772 483236
rect 573008 483092 573244 483328
rect 573480 483092 573716 483328
rect 573952 483092 574188 483328
rect 574424 483092 574660 483328
rect 574896 483092 575132 483328
rect 575368 483092 575604 483328
rect 575840 483092 576076 483328
rect 576312 483092 576548 483328
rect 576784 483092 577020 483328
rect 577256 483092 578504 483328
rect 536504 482856 578504 483092
rect 536504 482620 572772 482856
rect 573008 482620 573244 482856
rect 573480 482620 573716 482856
rect 573952 482620 574188 482856
rect 574424 482620 574660 482856
rect 574896 482620 575132 482856
rect 575368 482620 575604 482856
rect 575840 482620 576076 482856
rect 576312 482620 576548 482856
rect 576784 482620 577020 482856
rect 577256 482620 578504 482856
rect 536504 482384 578504 482620
rect 536504 482148 572772 482384
rect 573008 482148 573244 482384
rect 573480 482148 573716 482384
rect 573952 482148 574188 482384
rect 574424 482148 574660 482384
rect 574896 482148 575132 482384
rect 575368 482148 575604 482384
rect 575840 482148 576076 482384
rect 576312 482148 576548 482384
rect 576784 482148 577020 482384
rect 577256 482148 578504 482384
rect 536504 481912 578504 482148
rect 536504 481676 572772 481912
rect 573008 481676 573244 481912
rect 573480 481676 573716 481912
rect 573952 481676 574188 481912
rect 574424 481676 574660 481912
rect 574896 481676 575132 481912
rect 575368 481676 575604 481912
rect 575840 481676 576076 481912
rect 576312 481676 576548 481912
rect 576784 481676 577020 481912
rect 577256 481676 578504 481912
rect 536504 481440 578504 481676
rect 536504 481204 572772 481440
rect 573008 481204 573244 481440
rect 573480 481204 573716 481440
rect 573952 481204 574188 481440
rect 574424 481204 574660 481440
rect 574896 481204 575132 481440
rect 575368 481204 575604 481440
rect 575840 481204 576076 481440
rect 576312 481204 576548 481440
rect 576784 481204 577020 481440
rect 577256 481204 578504 481440
rect 536504 480968 578504 481204
rect 536504 480732 572772 480968
rect 573008 480732 573244 480968
rect 573480 480732 573716 480968
rect 573952 480732 574188 480968
rect 574424 480732 574660 480968
rect 574896 480732 575132 480968
rect 575368 480732 575604 480968
rect 575840 480732 576076 480968
rect 576312 480732 576548 480968
rect 576784 480732 577020 480968
rect 577256 480732 578504 480968
rect 536504 480496 578504 480732
rect 536504 480260 572772 480496
rect 573008 480260 573244 480496
rect 573480 480260 573716 480496
rect 573952 480260 574188 480496
rect 574424 480260 574660 480496
rect 574896 480260 575132 480496
rect 575368 480260 575604 480496
rect 575840 480260 576076 480496
rect 576312 480260 576548 480496
rect 576784 480260 577020 480496
rect 577256 480260 578504 480496
rect 536504 480024 578504 480260
rect 536504 479788 572772 480024
rect 573008 479788 573244 480024
rect 573480 479788 573716 480024
rect 573952 479788 574188 480024
rect 574424 479788 574660 480024
rect 574896 479788 575132 480024
rect 575368 479788 575604 480024
rect 575840 479788 576076 480024
rect 576312 479788 576548 480024
rect 576784 479788 577020 480024
rect 577256 479788 578504 480024
rect 536504 479552 578504 479788
rect 536504 479316 572772 479552
rect 573008 479316 573244 479552
rect 573480 479316 573716 479552
rect 573952 479316 574188 479552
rect 574424 479316 574660 479552
rect 574896 479316 575132 479552
rect 575368 479316 575604 479552
rect 575840 479316 576076 479552
rect 576312 479316 576548 479552
rect 576784 479316 577020 479552
rect 577256 479316 578504 479552
rect 536504 479080 578504 479316
rect 536504 478844 572772 479080
rect 573008 478844 573244 479080
rect 573480 478844 573716 479080
rect 573952 478844 574188 479080
rect 574424 478844 574660 479080
rect 574896 478844 575132 479080
rect 575368 478844 575604 479080
rect 575840 478844 576076 479080
rect 576312 478844 576548 479080
rect 576784 478844 577020 479080
rect 577256 478844 578504 479080
rect 536504 478608 578504 478844
rect 536504 478452 572772 478608
rect 490440 478372 572772 478452
rect 573008 478372 573244 478608
rect 573480 478372 573716 478608
rect 573952 478372 574188 478608
rect 574424 478372 574660 478608
rect 574896 478372 575132 478608
rect 575368 478372 575604 478608
rect 575840 478372 576076 478608
rect 576312 478372 576548 478608
rect 576784 478372 577020 478608
rect 577256 478372 578504 478608
rect 490440 478136 578504 478372
rect 490440 477900 572772 478136
rect 573008 477900 573244 478136
rect 573480 477900 573716 478136
rect 573952 477900 574188 478136
rect 574424 477900 574660 478136
rect 574896 477900 575132 478136
rect 575368 477900 575604 478136
rect 575840 477900 576076 478136
rect 576312 477900 576548 478136
rect 576784 477900 577020 478136
rect 577256 477900 578504 478136
rect 490440 477580 578504 477900
rect 503864 475336 510520 475436
rect 503864 475306 510526 475336
rect 503864 475206 503920 475306
rect 504020 475206 504144 475306
rect 504244 475206 504368 475306
rect 504468 475206 504592 475306
rect 504692 475206 504816 475306
rect 504916 475206 505040 475306
rect 505140 475206 505264 475306
rect 505364 475206 505488 475306
rect 505588 475206 505712 475306
rect 505812 475206 505936 475306
rect 506036 475206 506160 475306
rect 506260 475206 506384 475306
rect 506484 475206 506608 475306
rect 506708 475206 506832 475306
rect 506932 475206 507056 475306
rect 507156 475206 507280 475306
rect 507380 475206 507504 475306
rect 507604 475206 507728 475306
rect 507828 475206 507952 475306
rect 508052 475206 508176 475306
rect 508276 475206 508400 475306
rect 508500 475206 508624 475306
rect 508724 475206 508848 475306
rect 508948 475206 509072 475306
rect 509172 475206 509296 475306
rect 509396 475206 509520 475306
rect 509620 475206 509744 475306
rect 509844 475206 509968 475306
rect 510068 475206 510192 475306
rect 510292 475206 510416 475306
rect 510516 475206 510526 475306
rect 503864 475082 510526 475206
rect 503864 474982 503920 475082
rect 504020 474982 504144 475082
rect 504244 474982 504368 475082
rect 504468 474982 504592 475082
rect 504692 474982 504816 475082
rect 504916 474982 505040 475082
rect 505140 474982 505264 475082
rect 505364 474982 505488 475082
rect 505588 474982 505712 475082
rect 505812 474982 505936 475082
rect 506036 474982 506160 475082
rect 506260 474982 506384 475082
rect 506484 474982 506608 475082
rect 506708 474982 506832 475082
rect 506932 474982 507056 475082
rect 507156 474982 507280 475082
rect 507380 474982 507504 475082
rect 507604 474982 507728 475082
rect 507828 474982 507952 475082
rect 508052 474982 508176 475082
rect 508276 474982 508400 475082
rect 508500 474982 508624 475082
rect 508724 474982 508848 475082
rect 508948 474982 509072 475082
rect 509172 474982 509296 475082
rect 509396 474982 509520 475082
rect 509620 474982 509744 475082
rect 509844 474982 509968 475082
rect 510068 474982 510192 475082
rect 510292 474982 510416 475082
rect 510516 474982 510526 475082
rect 503864 474858 510526 474982
rect 503864 474758 503920 474858
rect 504020 474758 504144 474858
rect 504244 474758 504368 474858
rect 504468 474758 504592 474858
rect 504692 474758 504816 474858
rect 504916 474758 505040 474858
rect 505140 474758 505264 474858
rect 505364 474758 505488 474858
rect 505588 474758 505712 474858
rect 505812 474758 505936 474858
rect 506036 474758 506160 474858
rect 506260 474758 506384 474858
rect 506484 474758 506608 474858
rect 506708 474758 506832 474858
rect 506932 474758 507056 474858
rect 507156 474758 507280 474858
rect 507380 474758 507504 474858
rect 507604 474758 507728 474858
rect 507828 474758 507952 474858
rect 508052 474758 508176 474858
rect 508276 474758 508400 474858
rect 508500 474758 508624 474858
rect 508724 474758 508848 474858
rect 508948 474758 509072 474858
rect 509172 474758 509296 474858
rect 509396 474758 509520 474858
rect 509620 474758 509744 474858
rect 509844 474758 509968 474858
rect 510068 474758 510192 474858
rect 510292 474758 510416 474858
rect 510516 474758 510526 474858
rect 503864 474634 510526 474758
rect 503864 474534 503920 474634
rect 504020 474534 504144 474634
rect 504244 474534 504368 474634
rect 504468 474534 504592 474634
rect 504692 474534 504816 474634
rect 504916 474534 505040 474634
rect 505140 474534 505264 474634
rect 505364 474534 505488 474634
rect 505588 474534 505712 474634
rect 505812 474534 505936 474634
rect 506036 474534 506160 474634
rect 506260 474534 506384 474634
rect 506484 474534 506608 474634
rect 506708 474534 506832 474634
rect 506932 474534 507056 474634
rect 507156 474534 507280 474634
rect 507380 474534 507504 474634
rect 507604 474534 507728 474634
rect 507828 474534 507952 474634
rect 508052 474534 508176 474634
rect 508276 474534 508400 474634
rect 508500 474534 508624 474634
rect 508724 474534 508848 474634
rect 508948 474534 509072 474634
rect 509172 474534 509296 474634
rect 509396 474534 509520 474634
rect 509620 474534 509744 474634
rect 509844 474534 509968 474634
rect 510068 474534 510192 474634
rect 510292 474534 510416 474634
rect 510516 474534 510526 474634
rect 503864 474410 510526 474534
rect 490440 474280 501440 474336
rect 490440 474236 500398 474280
rect 490440 469452 491256 474236
rect 497000 474180 500398 474236
rect 500498 474180 500622 474280
rect 500722 474180 500846 474280
rect 500946 474180 501070 474280
rect 501170 474180 501294 474280
rect 501394 474180 501440 474280
rect 503864 474310 503920 474410
rect 504020 474310 504144 474410
rect 504244 474310 504368 474410
rect 504468 474310 504592 474410
rect 504692 474310 504816 474410
rect 504916 474310 505040 474410
rect 505140 474310 505264 474410
rect 505364 474310 505488 474410
rect 505588 474310 505712 474410
rect 505812 474310 505936 474410
rect 506036 474310 506160 474410
rect 506260 474310 506384 474410
rect 506484 474310 506608 474410
rect 506708 474310 506832 474410
rect 506932 474310 507056 474410
rect 507156 474310 507280 474410
rect 507380 474310 507504 474410
rect 507604 474310 507728 474410
rect 507828 474310 507952 474410
rect 508052 474310 508176 474410
rect 508276 474310 508400 474410
rect 508500 474310 508624 474410
rect 508724 474310 508848 474410
rect 508948 474310 509072 474410
rect 509172 474310 509296 474410
rect 509396 474310 509520 474410
rect 509620 474310 509744 474410
rect 509844 474310 509968 474410
rect 510068 474310 510192 474410
rect 510292 474310 510416 474410
rect 510516 474310 510526 474410
rect 503864 474278 510526 474310
rect 511584 475300 512160 475364
rect 511584 475236 511648 475300
rect 511712 475236 511776 475300
rect 511840 475236 511904 475300
rect 511968 475236 512032 475300
rect 512096 475236 512160 475300
rect 511584 475172 512160 475236
rect 511584 475108 511648 475172
rect 511712 475108 511776 475172
rect 511840 475108 511904 475172
rect 511968 475108 512032 475172
rect 512096 475108 512160 475172
rect 511584 475044 512160 475108
rect 511584 474980 511648 475044
rect 511712 474980 511776 475044
rect 511840 474980 511904 475044
rect 511968 474980 512032 475044
rect 512096 474980 512160 475044
rect 511584 474916 512160 474980
rect 511584 474852 511648 474916
rect 511712 474852 511776 474916
rect 511840 474852 511904 474916
rect 511968 474852 512032 474916
rect 512096 474852 512160 474916
rect 511584 474788 512160 474852
rect 511584 474724 511648 474788
rect 511712 474724 511776 474788
rect 511840 474724 511904 474788
rect 511968 474724 512032 474788
rect 512096 474724 512160 474788
rect 511584 474660 512160 474724
rect 511584 474596 511648 474660
rect 511712 474596 511776 474660
rect 511840 474596 511904 474660
rect 511968 474596 512032 474660
rect 512096 474596 512160 474660
rect 511584 474532 512160 474596
rect 511584 474468 511648 474532
rect 511712 474468 511776 474532
rect 511840 474468 511904 474532
rect 511968 474468 512032 474532
rect 512096 474468 512160 474532
rect 511584 474404 512160 474468
rect 511584 474340 511648 474404
rect 511712 474340 511776 474404
rect 511840 474340 511904 474404
rect 511968 474340 512032 474404
rect 512096 474340 512160 474404
rect 503864 474276 510520 474278
rect 511584 474276 512160 474340
rect 517280 475306 523940 475336
rect 517280 475206 517320 475306
rect 517420 475206 517544 475306
rect 517644 475206 517768 475306
rect 517868 475206 517992 475306
rect 518092 475206 518216 475306
rect 518316 475206 518440 475306
rect 518540 475206 518664 475306
rect 518764 475206 518888 475306
rect 518988 475206 519112 475306
rect 519212 475206 519336 475306
rect 519436 475206 519560 475306
rect 519660 475206 519784 475306
rect 519884 475206 520008 475306
rect 520108 475206 520232 475306
rect 520332 475206 520456 475306
rect 520556 475206 520680 475306
rect 520780 475206 520904 475306
rect 521004 475206 521128 475306
rect 521228 475206 521352 475306
rect 521452 475206 521576 475306
rect 521676 475206 521800 475306
rect 521900 475206 522024 475306
rect 522124 475206 522248 475306
rect 522348 475206 522472 475306
rect 522572 475206 522696 475306
rect 522796 475206 522920 475306
rect 523020 475206 523144 475306
rect 523244 475206 523368 475306
rect 523468 475206 523592 475306
rect 523692 475206 523816 475306
rect 523916 475206 523940 475306
rect 517280 475082 523940 475206
rect 517280 474982 517320 475082
rect 517420 474982 517544 475082
rect 517644 474982 517768 475082
rect 517868 474982 517992 475082
rect 518092 474982 518216 475082
rect 518316 474982 518440 475082
rect 518540 474982 518664 475082
rect 518764 474982 518888 475082
rect 518988 474982 519112 475082
rect 519212 474982 519336 475082
rect 519436 474982 519560 475082
rect 519660 474982 519784 475082
rect 519884 474982 520008 475082
rect 520108 474982 520232 475082
rect 520332 474982 520456 475082
rect 520556 474982 520680 475082
rect 520780 474982 520904 475082
rect 521004 474982 521128 475082
rect 521228 474982 521352 475082
rect 521452 474982 521576 475082
rect 521676 474982 521800 475082
rect 521900 474982 522024 475082
rect 522124 474982 522248 475082
rect 522348 474982 522472 475082
rect 522572 474982 522696 475082
rect 522796 474982 522920 475082
rect 523020 474982 523144 475082
rect 523244 474982 523368 475082
rect 523468 474982 523592 475082
rect 523692 474982 523816 475082
rect 523916 474982 523940 475082
rect 517280 474858 523940 474982
rect 517280 474758 517320 474858
rect 517420 474758 517544 474858
rect 517644 474758 517768 474858
rect 517868 474758 517992 474858
rect 518092 474758 518216 474858
rect 518316 474758 518440 474858
rect 518540 474758 518664 474858
rect 518764 474758 518888 474858
rect 518988 474758 519112 474858
rect 519212 474758 519336 474858
rect 519436 474758 519560 474858
rect 519660 474758 519784 474858
rect 519884 474758 520008 474858
rect 520108 474758 520232 474858
rect 520332 474758 520456 474858
rect 520556 474758 520680 474858
rect 520780 474758 520904 474858
rect 521004 474758 521128 474858
rect 521228 474758 521352 474858
rect 521452 474758 521576 474858
rect 521676 474758 521800 474858
rect 521900 474758 522024 474858
rect 522124 474758 522248 474858
rect 522348 474758 522472 474858
rect 522572 474758 522696 474858
rect 522796 474758 522920 474858
rect 523020 474758 523144 474858
rect 523244 474758 523368 474858
rect 523468 474758 523592 474858
rect 523692 474758 523816 474858
rect 523916 474758 523940 474858
rect 517280 474634 523940 474758
rect 517280 474534 517320 474634
rect 517420 474534 517544 474634
rect 517644 474534 517768 474634
rect 517868 474534 517992 474634
rect 518092 474534 518216 474634
rect 518316 474534 518440 474634
rect 518540 474534 518664 474634
rect 518764 474534 518888 474634
rect 518988 474534 519112 474634
rect 519212 474534 519336 474634
rect 519436 474534 519560 474634
rect 519660 474534 519784 474634
rect 519884 474534 520008 474634
rect 520108 474534 520232 474634
rect 520332 474534 520456 474634
rect 520556 474534 520680 474634
rect 520780 474534 520904 474634
rect 521004 474534 521128 474634
rect 521228 474534 521352 474634
rect 521452 474534 521576 474634
rect 521676 474534 521800 474634
rect 521900 474534 522024 474634
rect 522124 474534 522248 474634
rect 522348 474534 522472 474634
rect 522572 474534 522696 474634
rect 522796 474534 522920 474634
rect 523020 474534 523144 474634
rect 523244 474534 523368 474634
rect 523468 474534 523592 474634
rect 523692 474534 523816 474634
rect 523916 474534 523940 474634
rect 517280 474410 523940 474534
rect 517280 474310 517320 474410
rect 517420 474310 517544 474410
rect 517644 474310 517768 474410
rect 517868 474310 517992 474410
rect 518092 474310 518216 474410
rect 518316 474310 518440 474410
rect 518540 474310 518664 474410
rect 518764 474310 518888 474410
rect 518988 474310 519112 474410
rect 519212 474310 519336 474410
rect 519436 474310 519560 474410
rect 519660 474310 519784 474410
rect 519884 474310 520008 474410
rect 520108 474310 520232 474410
rect 520332 474310 520456 474410
rect 520556 474310 520680 474410
rect 520780 474310 520904 474410
rect 521004 474310 521128 474410
rect 521228 474310 521352 474410
rect 521452 474310 521576 474410
rect 521676 474310 521800 474410
rect 521900 474310 522024 474410
rect 522124 474310 522248 474410
rect 522348 474310 522472 474410
rect 522572 474310 522696 474410
rect 522796 474310 522920 474410
rect 523020 474310 523144 474410
rect 523244 474310 523368 474410
rect 523468 474310 523592 474410
rect 523692 474310 523816 474410
rect 523916 474310 523940 474410
rect 517280 474276 523940 474310
rect 527580 474280 537320 474336
rect 497000 474056 501440 474180
rect 497000 473956 500398 474056
rect 500498 473956 500622 474056
rect 500722 473956 500846 474056
rect 500946 473956 501070 474056
rect 501170 473956 501294 474056
rect 501394 473956 501440 474056
rect 497000 473832 501440 473956
rect 497000 473732 500398 473832
rect 500498 473732 500622 473832
rect 500722 473732 500846 473832
rect 500946 473732 501070 473832
rect 501170 473732 501294 473832
rect 501394 473732 501440 473832
rect 497000 473608 501440 473732
rect 497000 473508 500398 473608
rect 500498 473508 500622 473608
rect 500722 473508 500846 473608
rect 500946 473508 501070 473608
rect 501170 473508 501294 473608
rect 501394 473508 501440 473608
rect 497000 473384 501440 473508
rect 497000 473284 500398 473384
rect 500498 473284 500622 473384
rect 500722 473284 500846 473384
rect 500946 473284 501070 473384
rect 501170 473284 501294 473384
rect 501394 473284 501440 473384
rect 497000 473160 501440 473284
rect 497000 473060 500398 473160
rect 500498 473060 500622 473160
rect 500722 473060 500846 473160
rect 500946 473060 501070 473160
rect 501170 473060 501294 473160
rect 501394 473060 501440 473160
rect 497000 472936 501440 473060
rect 497000 472836 500398 472936
rect 500498 472836 500622 472936
rect 500722 472836 500846 472936
rect 500946 472836 501070 472936
rect 501170 472836 501294 472936
rect 501394 472836 501440 472936
rect 497000 472712 501440 472836
rect 497000 472612 500398 472712
rect 500498 472612 500622 472712
rect 500722 472612 500846 472712
rect 500946 472612 501070 472712
rect 501170 472612 501294 472712
rect 501394 472612 501440 472712
rect 497000 472488 501440 472612
rect 497000 472388 500398 472488
rect 500498 472388 500622 472488
rect 500722 472388 500846 472488
rect 500946 472388 501070 472488
rect 501170 472388 501294 472488
rect 501394 472388 501440 472488
rect 497000 472264 501440 472388
rect 497000 472164 500398 472264
rect 500498 472164 500622 472264
rect 500722 472164 500846 472264
rect 500946 472164 501070 472264
rect 501170 472164 501294 472264
rect 501394 472164 501440 472264
rect 497000 472040 501440 472164
rect 497000 471940 500398 472040
rect 500498 471940 500622 472040
rect 500722 471940 500846 472040
rect 500946 471940 501070 472040
rect 501170 471940 501294 472040
rect 501394 471940 501440 472040
rect 497000 471816 501440 471940
rect 497000 471716 500398 471816
rect 500498 471716 500622 471816
rect 500722 471716 500846 471816
rect 500946 471716 501070 471816
rect 501170 471716 501294 471816
rect 501394 471716 501440 471816
rect 497000 471592 501440 471716
rect 497000 471492 500398 471592
rect 500498 471492 500622 471592
rect 500722 471492 500846 471592
rect 500946 471492 501070 471592
rect 501170 471492 501294 471592
rect 501394 471492 501440 471592
rect 497000 471368 501440 471492
rect 497000 471268 500398 471368
rect 500498 471268 500622 471368
rect 500722 471268 500846 471368
rect 500946 471268 501070 471368
rect 501170 471268 501294 471368
rect 501394 471268 501440 471368
rect 497000 471144 501440 471268
rect 511584 474212 511648 474276
rect 511712 474212 511776 474276
rect 511840 474212 511904 474276
rect 511968 474212 512032 474276
rect 512096 474212 512160 474276
rect 497000 471044 500398 471144
rect 500498 471044 500622 471144
rect 500722 471044 500846 471144
rect 500946 471044 501070 471144
rect 501170 471044 501294 471144
rect 501394 471044 501440 471144
rect 497000 470920 501440 471044
rect 497000 470820 500398 470920
rect 500498 470820 500622 470920
rect 500722 470820 500846 470920
rect 500946 470820 501070 470920
rect 501170 470820 501294 470920
rect 501394 470820 501440 470920
rect 497000 470696 501440 470820
rect 497000 470596 500398 470696
rect 500498 470596 500622 470696
rect 500722 470596 500846 470696
rect 500946 470596 501070 470696
rect 501170 470596 501294 470696
rect 501394 470596 501440 470696
rect 497000 470472 501440 470596
rect 497000 470372 500398 470472
rect 500498 470372 500622 470472
rect 500722 470372 500846 470472
rect 500946 470372 501070 470472
rect 501170 470372 501294 470472
rect 501394 470372 501440 470472
rect 497000 470248 501440 470372
rect 497000 470148 500398 470248
rect 500498 470148 500622 470248
rect 500722 470148 500846 470248
rect 500946 470148 501070 470248
rect 501170 470148 501294 470248
rect 501394 470148 501440 470248
rect 497000 470024 501440 470148
rect 497000 469924 500398 470024
rect 500498 469924 500622 470024
rect 500722 469924 500846 470024
rect 500946 469924 501070 470024
rect 501170 469924 501294 470024
rect 501394 469924 501440 470024
rect 497000 469800 501440 469924
rect 497000 469700 500398 469800
rect 500498 469700 500622 469800
rect 500722 469700 500846 469800
rect 500946 469700 501070 469800
rect 501170 469700 501294 469800
rect 501394 469700 501440 469800
rect 497000 469576 501440 469700
rect 497000 469476 500398 469576
rect 500498 469476 500622 469576
rect 500722 469476 500846 469576
rect 500946 469476 501070 469576
rect 501170 469476 501294 469576
rect 501394 469476 501440 469576
rect 497000 469452 501440 469476
rect 490440 469352 501440 469452
rect 490440 469252 500398 469352
rect 500498 469252 500622 469352
rect 500722 469252 500846 469352
rect 500946 469252 501070 469352
rect 501170 469252 501294 469352
rect 501394 469252 501440 469352
rect 490440 469128 501440 469252
rect 490440 469028 500398 469128
rect 500498 469028 500622 469128
rect 500722 469028 500846 469128
rect 500946 469028 501070 469128
rect 501170 469028 501294 469128
rect 501394 469028 501440 469128
rect 490440 468904 501440 469028
rect 490440 468804 500398 468904
rect 500498 468804 500622 468904
rect 500722 468804 500846 468904
rect 500946 468804 501070 468904
rect 501170 468804 501294 468904
rect 501394 468804 501440 468904
rect 502426 470218 502868 471218
rect 502426 470210 502988 470218
rect 502426 468840 502868 470210
rect 490440 468680 501440 468804
rect 490440 468580 500398 468680
rect 500498 468580 500622 468680
rect 500722 468580 500846 468680
rect 500946 468580 501070 468680
rect 501170 468580 501294 468680
rect 501394 468580 501440 468680
rect 490440 468456 501440 468580
rect -800 468308 480 468420
rect 490440 468356 500398 468456
rect 500498 468356 500622 468456
rect 500722 468356 500846 468456
rect 500946 468356 501070 468456
rect 501170 468356 501294 468456
rect 501394 468356 501440 468456
rect 490440 468236 501440 468356
rect -800 467126 480 467238
rect -800 465944 480 466056
rect -800 464762 480 464874
rect -800 463580 480 463692
rect 490440 463452 491256 468236
rect 497000 468232 501440 468236
rect 497000 468132 500398 468232
rect 500498 468132 500622 468232
rect 500722 468132 500846 468232
rect 500946 468132 501070 468232
rect 501170 468132 501294 468232
rect 501394 468132 501440 468232
rect 497000 468008 501440 468132
rect 497000 467908 500398 468008
rect 500498 467908 500622 468008
rect 500722 467908 500846 468008
rect 500946 467908 501070 468008
rect 501170 467908 501294 468008
rect 501394 467908 501440 468008
rect 497000 467784 501440 467908
rect 497000 467684 500398 467784
rect 500498 467684 500622 467784
rect 500722 467684 500846 467784
rect 500946 467684 501070 467784
rect 501170 467684 501294 467784
rect 501394 467684 501440 467784
rect 497000 463810 501440 467684
rect 497000 463710 500398 463810
rect 500498 463710 500622 463810
rect 500722 463710 500846 463810
rect 500946 463710 501070 463810
rect 501170 463710 501294 463810
rect 501394 463710 501440 463810
rect 497000 463586 501440 463710
rect 497000 463486 500398 463586
rect 500498 463486 500622 463586
rect 500722 463486 500846 463586
rect 500946 463486 501070 463586
rect 501170 463486 501294 463586
rect 501394 463486 501440 463586
rect 497000 463452 501440 463486
rect 490440 463362 501440 463452
rect 490440 463262 500398 463362
rect 500498 463262 500622 463362
rect 500722 463262 500846 463362
rect 500946 463262 501070 463362
rect 501170 463262 501294 463362
rect 501394 463262 501440 463362
rect 490440 463138 501440 463262
rect 490440 463038 500398 463138
rect 500498 463038 500622 463138
rect 500722 463038 500846 463138
rect 500946 463038 501070 463138
rect 501170 463038 501294 463138
rect 501394 463038 501440 463138
rect 490440 462914 501440 463038
rect 490440 462814 500398 462914
rect 500498 462814 500622 462914
rect 500722 462814 500846 462914
rect 500946 462814 501070 462914
rect 501170 462814 501294 462914
rect 501394 462814 501440 462914
rect 490440 462690 501440 462814
rect 490440 462590 500398 462690
rect 500498 462590 500622 462690
rect 500722 462590 500846 462690
rect 500946 462590 501070 462690
rect 501170 462590 501294 462690
rect 501394 462590 501440 462690
rect -800 462398 480 462510
rect 490440 462466 501440 462590
rect 490440 462366 500398 462466
rect 500498 462366 500622 462466
rect 500722 462366 500846 462466
rect 500946 462366 501070 462466
rect 501170 462366 501294 462466
rect 501394 462366 501440 462466
rect 490440 462242 501440 462366
rect 490440 462236 500398 462242
rect 490440 457452 491256 462236
rect 497000 462142 500398 462236
rect 500498 462142 500622 462242
rect 500722 462142 500846 462242
rect 500946 462142 501070 462242
rect 501170 462142 501294 462242
rect 501394 462142 501440 462242
rect 497000 462018 501440 462142
rect 497000 461918 500398 462018
rect 500498 461918 500622 462018
rect 500722 461918 500846 462018
rect 500946 461918 501070 462018
rect 501170 461918 501294 462018
rect 501394 461918 501440 462018
rect 497000 461794 501440 461918
rect 497000 461694 500398 461794
rect 500498 461694 500622 461794
rect 500722 461694 500846 461794
rect 500946 461694 501070 461794
rect 501170 461694 501294 461794
rect 501394 461694 501440 461794
rect 497000 461570 501440 461694
rect 502392 461670 502868 468840
rect 497000 461470 500398 461570
rect 500498 461470 500622 461570
rect 500722 461470 500846 461570
rect 500946 461470 501070 461570
rect 501170 461470 501294 461570
rect 501394 461470 501440 461570
rect 497000 461346 501440 461470
rect 497000 461246 500398 461346
rect 500498 461246 500622 461346
rect 500722 461246 500846 461346
rect 500946 461246 501070 461346
rect 501170 461246 501294 461346
rect 501394 461246 501440 461346
rect 497000 461122 501440 461246
rect 497000 461022 500398 461122
rect 500498 461022 500622 461122
rect 500722 461022 500846 461122
rect 500946 461022 501070 461122
rect 501170 461022 501294 461122
rect 501394 461022 501440 461122
rect 497000 460898 501440 461022
rect 497000 460798 500398 460898
rect 500498 460798 500622 460898
rect 500722 460798 500846 460898
rect 500946 460798 501070 460898
rect 501170 460798 501294 460898
rect 501394 460798 501440 460898
rect 497000 460674 501440 460798
rect 497000 460574 500398 460674
rect 500498 460574 500622 460674
rect 500722 460574 500846 460674
rect 500946 460574 501070 460674
rect 501170 460574 501294 460674
rect 501394 460574 501440 460674
rect 497000 460450 501440 460574
rect 497000 460350 500398 460450
rect 500498 460350 500622 460450
rect 500722 460350 500846 460450
rect 500946 460350 501070 460450
rect 501170 460350 501294 460450
rect 501394 460350 501440 460450
rect 497000 460226 501440 460350
rect 497000 460126 500398 460226
rect 500498 460126 500622 460226
rect 500722 460126 500846 460226
rect 500946 460126 501070 460226
rect 501170 460126 501294 460226
rect 501394 460126 501440 460226
rect 497000 460002 501440 460126
rect 497000 459902 500398 460002
rect 500498 459902 500622 460002
rect 500722 459902 500846 460002
rect 500946 459902 501070 460002
rect 501170 459902 501294 460002
rect 501394 459902 501440 460002
rect 497000 459778 501440 459902
rect 497000 459678 500398 459778
rect 500498 459678 500622 459778
rect 500722 459678 500846 459778
rect 500946 459678 501070 459778
rect 501170 459678 501294 459778
rect 501394 459678 501440 459778
rect 497000 459554 501440 459678
rect 497000 459454 500398 459554
rect 500498 459454 500622 459554
rect 500722 459454 500846 459554
rect 500946 459454 501070 459554
rect 501170 459454 501294 459554
rect 501394 459454 501440 459554
rect 497000 459330 501440 459454
rect 497000 459230 500398 459330
rect 500498 459230 500622 459330
rect 500722 459230 500846 459330
rect 500946 459230 501070 459330
rect 501170 459230 501294 459330
rect 501394 459230 501440 459330
rect 497000 459106 501440 459230
rect 497000 459006 500398 459106
rect 500498 459006 500622 459106
rect 500722 459006 500846 459106
rect 500946 459006 501070 459106
rect 501170 459006 501294 459106
rect 501394 459006 501440 459106
rect 497000 458882 501440 459006
rect 497000 458782 500398 458882
rect 500498 458782 500622 458882
rect 500722 458782 500846 458882
rect 500946 458782 501070 458882
rect 501170 458782 501294 458882
rect 501394 458782 501440 458882
rect 497000 458658 501440 458782
rect 497000 458558 500398 458658
rect 500498 458558 500622 458658
rect 500722 458558 500846 458658
rect 500946 458558 501070 458658
rect 501170 458558 501294 458658
rect 501394 458558 501440 458658
rect 497000 458434 501440 458558
rect 497000 458334 500398 458434
rect 500498 458334 500622 458434
rect 500722 458334 500846 458434
rect 500946 458334 501070 458434
rect 501170 458334 501294 458434
rect 501394 458334 501440 458434
rect 497000 458210 501440 458334
rect 497000 458110 500398 458210
rect 500498 458110 500622 458210
rect 500722 458110 500846 458210
rect 500946 458110 501070 458210
rect 501170 458110 501294 458210
rect 501394 458110 501440 458210
rect 497000 457986 501440 458110
rect 497000 457886 500398 457986
rect 500498 457886 500622 457986
rect 500722 457886 500846 457986
rect 500946 457886 501070 457986
rect 501170 457886 501294 457986
rect 501394 457886 501440 457986
rect 497000 457762 501440 457886
rect 497000 457662 500398 457762
rect 500498 457662 500622 457762
rect 500722 457662 500846 457762
rect 500946 457662 501070 457762
rect 501170 457662 501294 457762
rect 501394 457662 501440 457762
rect 497000 457538 501440 457662
rect 497000 457452 500398 457538
rect 490440 457438 500398 457452
rect 500498 457438 500622 457538
rect 500722 457438 500846 457538
rect 500946 457438 501070 457538
rect 501170 457438 501294 457538
rect 501394 457438 501440 457538
rect 490440 457314 501440 457438
rect 490440 457214 500398 457314
rect 500498 457214 500622 457314
rect 500722 457214 500846 457314
rect 500946 457214 501070 457314
rect 501170 457214 501294 457314
rect 501394 457214 501440 457314
rect 490440 457196 501440 457214
rect 502426 460964 502868 461670
rect 502982 468840 502988 470210
rect 511584 470176 512160 474212
rect 527580 474180 527618 474280
rect 527718 474180 527842 474280
rect 527942 474180 528066 474280
rect 528166 474180 528290 474280
rect 528390 474180 528514 474280
rect 528614 474236 537320 474280
rect 528614 474180 530760 474236
rect 527580 474056 530760 474180
rect 527580 473956 527618 474056
rect 527718 473956 527842 474056
rect 527942 473956 528066 474056
rect 528166 473956 528290 474056
rect 528390 473956 528514 474056
rect 528614 473956 530760 474056
rect 527580 473832 530760 473956
rect 527580 473732 527618 473832
rect 527718 473732 527842 473832
rect 527942 473732 528066 473832
rect 528166 473732 528290 473832
rect 528390 473732 528514 473832
rect 528614 473732 530760 473832
rect 527580 473608 530760 473732
rect 527580 473508 527618 473608
rect 527718 473508 527842 473608
rect 527942 473508 528066 473608
rect 528166 473508 528290 473608
rect 528390 473508 528514 473608
rect 528614 473508 530760 473608
rect 527580 473384 530760 473508
rect 527580 473284 527618 473384
rect 527718 473284 527842 473384
rect 527942 473284 528066 473384
rect 528166 473284 528290 473384
rect 528390 473284 528514 473384
rect 528614 473284 530760 473384
rect 527580 473160 530760 473284
rect 527580 473060 527618 473160
rect 527718 473060 527842 473160
rect 527942 473060 528066 473160
rect 528166 473060 528290 473160
rect 528390 473060 528514 473160
rect 528614 473060 530760 473160
rect 527580 472936 530760 473060
rect 527580 472836 527618 472936
rect 527718 472836 527842 472936
rect 527942 472836 528066 472936
rect 528166 472836 528290 472936
rect 528390 472836 528514 472936
rect 528614 472836 530760 472936
rect 527580 472712 530760 472836
rect 527580 472612 527618 472712
rect 527718 472612 527842 472712
rect 527942 472612 528066 472712
rect 528166 472612 528290 472712
rect 528390 472612 528514 472712
rect 528614 472612 530760 472712
rect 511584 470116 511770 470176
rect 511830 470116 511890 470176
rect 511950 470116 512160 470176
rect 511584 470056 512160 470116
rect 511584 469996 511770 470056
rect 511830 469996 511890 470056
rect 511950 469996 512160 470056
rect 511584 469936 512160 469996
rect 511584 469876 511770 469936
rect 511830 469876 511890 469936
rect 511950 469876 512160 469936
rect 511584 469816 512160 469876
rect 511584 469756 511770 469816
rect 511830 469756 511890 469816
rect 511950 469756 512160 469816
rect 511584 469696 512160 469756
rect 511584 469636 511770 469696
rect 511830 469636 511890 469696
rect 511950 469636 512160 469696
rect 511584 469604 512160 469636
rect 525645 472513 526513 472519
rect 505783 469566 506075 469572
rect 505783 468938 505789 469566
rect 506069 468938 506075 469566
rect 505783 468932 506075 468938
rect 502982 468225 518092 468840
rect 502982 468161 511220 468225
rect 511764 468161 511920 468225
rect 512464 468161 512620 468225
rect 513164 468161 513320 468225
rect 513864 468161 514020 468225
rect 514564 468161 514720 468225
rect 515264 468161 515420 468225
rect 515964 468161 516120 468225
rect 516664 468161 516820 468225
rect 517364 468161 517520 468225
rect 518064 468161 518092 468225
rect 502982 467506 518092 468161
rect 502982 467442 511220 467506
rect 511764 467442 511920 467506
rect 512464 467442 512620 467506
rect 513164 467442 513320 467506
rect 513864 467442 514020 467506
rect 514564 467442 514720 467506
rect 515264 467442 515420 467506
rect 515964 467442 516120 467506
rect 516664 467442 516820 467506
rect 517364 467442 517520 467506
rect 518064 467442 518092 467506
rect 502982 466787 518092 467442
rect 502982 466723 511220 466787
rect 511764 466723 511920 466787
rect 512464 466723 512620 466787
rect 513164 466723 513320 466787
rect 513864 466723 514020 466787
rect 514564 466723 514720 466787
rect 515264 466723 515420 466787
rect 515964 466723 516120 466787
rect 516664 466723 516820 466787
rect 517364 466723 517520 466787
rect 518064 466723 518092 466787
rect 502982 466068 518092 466723
rect 502982 466004 511220 466068
rect 511764 466004 511920 466068
rect 512464 466004 512620 466068
rect 513164 466004 513320 466068
rect 513864 466004 514020 466068
rect 514564 466004 514720 466068
rect 515264 466004 515420 466068
rect 515964 466004 516120 466068
rect 516664 466004 516820 466068
rect 517364 466004 517520 466068
rect 518064 466004 518092 466068
rect 502982 465349 518092 466004
rect 502982 465285 511220 465349
rect 511764 465285 511920 465349
rect 512464 465285 512620 465349
rect 513164 465285 513320 465349
rect 513864 465285 514020 465349
rect 514564 465285 514720 465349
rect 515264 465285 515420 465349
rect 515964 465285 516120 465349
rect 516664 465285 516820 465349
rect 517364 465285 517520 465349
rect 518064 465285 518092 465349
rect 502982 464630 518092 465285
rect 502982 464566 511220 464630
rect 511764 464566 511920 464630
rect 512464 464566 512620 464630
rect 513164 464566 513320 464630
rect 513864 464566 514020 464630
rect 514564 464566 514720 464630
rect 515264 464566 515420 464630
rect 515964 464566 516120 464630
rect 516664 464566 516820 464630
rect 517364 464566 517520 464630
rect 518064 464566 518092 464630
rect 502982 463911 518092 464566
rect 502982 463847 511220 463911
rect 511764 463847 511920 463911
rect 512464 463847 512620 463911
rect 513164 463847 513320 463911
rect 513864 463847 514020 463911
rect 514564 463847 514720 463911
rect 515264 463847 515420 463911
rect 515964 463847 516120 463911
rect 516664 463847 516820 463911
rect 517364 463847 517520 463911
rect 518064 463847 518092 463911
rect 502982 463192 518092 463847
rect 502982 463128 511220 463192
rect 511764 463128 511920 463192
rect 512464 463128 512620 463192
rect 513164 463128 513320 463192
rect 513864 463128 514020 463192
rect 514564 463128 514720 463192
rect 515264 463128 515420 463192
rect 515964 463128 516120 463192
rect 516664 463128 516820 463192
rect 517364 463128 517520 463192
rect 518064 463128 518092 463192
rect 502982 462473 518092 463128
rect 502982 462409 511220 462473
rect 511764 462409 511920 462473
rect 512464 462409 512620 462473
rect 513164 462409 513320 462473
rect 513864 462409 514020 462473
rect 514564 462409 514720 462473
rect 515264 462409 515420 462473
rect 515964 462409 516120 462473
rect 516664 462409 516820 462473
rect 517364 462409 517520 462473
rect 518064 462409 518092 462473
rect 502982 461754 518092 462409
rect 502982 461690 511220 461754
rect 511764 461690 511920 461754
rect 512464 461690 512620 461754
rect 513164 461690 513320 461754
rect 513864 461690 514020 461754
rect 514564 461690 514720 461754
rect 515264 461690 515420 461754
rect 515964 461690 516120 461754
rect 516664 461690 516820 461754
rect 517364 461690 517520 461754
rect 518064 461690 518092 461754
rect 502982 461670 518092 461690
rect 502982 460964 502988 461670
rect 525645 461239 525651 472513
rect 526507 461239 526513 472513
rect 525645 461233 526513 461239
rect 527580 472488 530760 472612
rect 527580 472388 527618 472488
rect 527718 472388 527842 472488
rect 527942 472388 528066 472488
rect 528166 472388 528290 472488
rect 528390 472388 528514 472488
rect 528614 472388 530760 472488
rect 527580 472264 530760 472388
rect 527580 472164 527618 472264
rect 527718 472164 527842 472264
rect 527942 472164 528066 472264
rect 528166 472164 528290 472264
rect 528390 472164 528514 472264
rect 528614 472164 530760 472264
rect 527580 472040 530760 472164
rect 527580 471940 527618 472040
rect 527718 471940 527842 472040
rect 527942 471940 528066 472040
rect 528166 471940 528290 472040
rect 528390 471940 528514 472040
rect 528614 471940 530760 472040
rect 527580 471816 530760 471940
rect 527580 471716 527618 471816
rect 527718 471716 527842 471816
rect 527942 471716 528066 471816
rect 528166 471716 528290 471816
rect 528390 471716 528514 471816
rect 528614 471716 530760 471816
rect 527580 471592 530760 471716
rect 527580 471492 527618 471592
rect 527718 471492 527842 471592
rect 527942 471492 528066 471592
rect 528166 471492 528290 471592
rect 528390 471492 528514 471592
rect 528614 471492 530760 471592
rect 527580 471368 530760 471492
rect 527580 471268 527618 471368
rect 527718 471268 527842 471368
rect 527942 471268 528066 471368
rect 528166 471268 528290 471368
rect 528390 471268 528514 471368
rect 528614 471268 530760 471368
rect 527580 471144 530760 471268
rect 527580 471044 527618 471144
rect 527718 471044 527842 471144
rect 527942 471044 528066 471144
rect 528166 471044 528290 471144
rect 528390 471044 528514 471144
rect 528614 471044 530760 471144
rect 527580 470920 530760 471044
rect 527580 470820 527618 470920
rect 527718 470820 527842 470920
rect 527942 470820 528066 470920
rect 528166 470820 528290 470920
rect 528390 470820 528514 470920
rect 528614 470820 530760 470920
rect 527580 470696 530760 470820
rect 527580 470596 527618 470696
rect 527718 470596 527842 470696
rect 527942 470596 528066 470696
rect 528166 470596 528290 470696
rect 528390 470596 528514 470696
rect 528614 470596 530760 470696
rect 527580 470472 530760 470596
rect 527580 470372 527618 470472
rect 527718 470372 527842 470472
rect 527942 470372 528066 470472
rect 528166 470372 528290 470472
rect 528390 470372 528514 470472
rect 528614 470372 530760 470472
rect 527580 470248 530760 470372
rect 527580 470148 527618 470248
rect 527718 470148 527842 470248
rect 527942 470148 528066 470248
rect 528166 470148 528290 470248
rect 528390 470148 528514 470248
rect 528614 470148 530760 470248
rect 527580 470024 530760 470148
rect 527580 469924 527618 470024
rect 527718 469924 527842 470024
rect 527942 469924 528066 470024
rect 528166 469924 528290 470024
rect 528390 469924 528514 470024
rect 528614 469924 530760 470024
rect 527580 469800 530760 469924
rect 527580 469700 527618 469800
rect 527718 469700 527842 469800
rect 527942 469700 528066 469800
rect 528166 469700 528290 469800
rect 528390 469700 528514 469800
rect 528614 469700 530760 469800
rect 527580 469576 530760 469700
rect 527580 469476 527618 469576
rect 527718 469476 527842 469576
rect 527942 469476 528066 469576
rect 528166 469476 528290 469576
rect 528390 469476 528514 469576
rect 528614 469476 530760 469576
rect 527580 469452 530760 469476
rect 536504 469452 537320 474236
rect 527580 469352 537320 469452
rect 527580 469252 527618 469352
rect 527718 469252 527842 469352
rect 527942 469252 528066 469352
rect 528166 469252 528290 469352
rect 528390 469252 528514 469352
rect 528614 469252 537320 469352
rect 527580 469128 537320 469252
rect 527580 469028 527618 469128
rect 527718 469028 527842 469128
rect 527942 469028 528066 469128
rect 528166 469028 528290 469128
rect 528390 469028 528514 469128
rect 528614 469028 537320 469128
rect 527580 468904 537320 469028
rect 527580 468804 527618 468904
rect 527718 468804 527842 468904
rect 527942 468804 528066 468904
rect 528166 468804 528290 468904
rect 528390 468804 528514 468904
rect 528614 468804 537320 468904
rect 527580 468680 537320 468804
rect 527580 468580 527618 468680
rect 527718 468580 527842 468680
rect 527942 468580 528066 468680
rect 528166 468580 528290 468680
rect 528390 468580 528514 468680
rect 528614 468580 537320 468680
rect 527580 468456 537320 468580
rect 527580 468356 527618 468456
rect 527718 468356 527842 468456
rect 527942 468356 528066 468456
rect 528166 468356 528290 468456
rect 528390 468356 528514 468456
rect 528614 468356 537320 468456
rect 527580 468236 537320 468356
rect 527580 468232 530760 468236
rect 527580 468132 527618 468232
rect 527718 468132 527842 468232
rect 527942 468132 528066 468232
rect 528166 468132 528290 468232
rect 528390 468132 528514 468232
rect 528614 468132 530760 468232
rect 527580 468008 530760 468132
rect 527580 467908 527618 468008
rect 527718 467908 527842 468008
rect 527942 467908 528066 468008
rect 528166 467908 528290 468008
rect 528390 467908 528514 468008
rect 528614 467908 530760 468008
rect 527580 467784 530760 467908
rect 527580 467684 527618 467784
rect 527718 467684 527842 467784
rect 527942 467684 528066 467784
rect 528166 467684 528290 467784
rect 528390 467684 528514 467784
rect 528614 467684 530760 467784
rect 527580 463810 530760 467684
rect 527580 463710 527618 463810
rect 527718 463710 527842 463810
rect 527942 463710 528066 463810
rect 528166 463710 528290 463810
rect 528390 463710 528514 463810
rect 528614 463710 530760 463810
rect 527580 463586 530760 463710
rect 527580 463486 527618 463586
rect 527718 463486 527842 463586
rect 527942 463486 528066 463586
rect 528166 463486 528290 463586
rect 528390 463486 528514 463586
rect 528614 463486 530760 463586
rect 527580 463452 530760 463486
rect 536504 463452 537320 468236
rect 527580 463362 537320 463452
rect 527580 463262 527618 463362
rect 527718 463262 527842 463362
rect 527942 463262 528066 463362
rect 528166 463262 528290 463362
rect 528390 463262 528514 463362
rect 528614 463262 537320 463362
rect 527580 463138 537320 463262
rect 527580 463038 527618 463138
rect 527718 463038 527842 463138
rect 527942 463038 528066 463138
rect 528166 463038 528290 463138
rect 528390 463038 528514 463138
rect 528614 463038 537320 463138
rect 527580 462914 537320 463038
rect 527580 462814 527618 462914
rect 527718 462814 527842 462914
rect 527942 462814 528066 462914
rect 528166 462814 528290 462914
rect 528390 462814 528514 462914
rect 528614 462814 537320 462914
rect 527580 462690 537320 462814
rect 527580 462590 527618 462690
rect 527718 462590 527842 462690
rect 527942 462590 528066 462690
rect 528166 462590 528290 462690
rect 528390 462590 528514 462690
rect 528614 462590 537320 462690
rect 527580 462466 537320 462590
rect 527580 462366 527618 462466
rect 527718 462366 527842 462466
rect 527942 462366 528066 462466
rect 528166 462366 528290 462466
rect 528390 462366 528514 462466
rect 528614 462366 537320 462466
rect 527580 462242 537320 462366
rect 527580 462142 527618 462242
rect 527718 462142 527842 462242
rect 527942 462142 528066 462242
rect 528166 462142 528290 462242
rect 528390 462142 528514 462242
rect 528614 462236 537320 462242
rect 528614 462142 530760 462236
rect 527580 462018 530760 462142
rect 527580 461918 527618 462018
rect 527718 461918 527842 462018
rect 527942 461918 528066 462018
rect 528166 461918 528290 462018
rect 528390 461918 528514 462018
rect 528614 461918 530760 462018
rect 527580 461794 530760 461918
rect 527580 461694 527618 461794
rect 527718 461694 527842 461794
rect 527942 461694 528066 461794
rect 528166 461694 528290 461794
rect 528390 461694 528514 461794
rect 528614 461694 530760 461794
rect 527580 461570 530760 461694
rect 527580 461470 527618 461570
rect 527718 461470 527842 461570
rect 527942 461470 528066 461570
rect 528166 461470 528290 461570
rect 528390 461470 528514 461570
rect 528614 461470 530760 461570
rect 527580 461346 530760 461470
rect 527580 461246 527618 461346
rect 527718 461246 527842 461346
rect 527942 461246 528066 461346
rect 528166 461246 528290 461346
rect 528390 461246 528514 461346
rect 528614 461246 530760 461346
rect 527580 461122 530760 461246
rect 502426 460446 502988 460964
rect 490440 457176 499020 457196
rect 502426 456196 502432 460446
rect 477000 455676 502432 456196
rect 477000 450892 477500 455676
rect 483244 450892 502432 455676
rect 477000 447676 502432 450892
rect 477000 442892 477500 447676
rect 483244 442892 502432 447676
rect 477000 442508 502432 442892
rect 502750 442508 502988 460446
rect 505783 461075 506075 461081
rect 505783 460447 505789 461075
rect 506069 460447 506075 461075
rect 505783 460441 506075 460447
rect 527580 461022 527618 461122
rect 527718 461022 527842 461122
rect 527942 461022 528066 461122
rect 528166 461022 528290 461122
rect 528390 461022 528514 461122
rect 528614 461022 530760 461122
rect 527580 460898 530760 461022
rect 527580 460798 527618 460898
rect 527718 460798 527842 460898
rect 527942 460798 528066 460898
rect 528166 460798 528290 460898
rect 528390 460798 528514 460898
rect 528614 460798 530760 460898
rect 527580 460674 530760 460798
rect 527580 460574 527618 460674
rect 527718 460574 527842 460674
rect 527942 460574 528066 460674
rect 528166 460574 528290 460674
rect 528390 460574 528514 460674
rect 528614 460574 530760 460674
rect 527580 460450 530760 460574
rect 527580 460350 527618 460450
rect 527718 460350 527842 460450
rect 527942 460350 528066 460450
rect 528166 460350 528290 460450
rect 528390 460350 528514 460450
rect 528614 460350 530760 460450
rect 527580 460226 530760 460350
rect 477000 442487 502988 442508
rect 512223 460204 513217 460209
rect 477000 442486 502766 442487
rect 477000 442476 502760 442486
rect 512223 439882 512228 460204
rect 513212 439882 513217 460204
rect 527580 460126 527618 460226
rect 527718 460126 527842 460226
rect 527942 460126 528066 460226
rect 528166 460126 528290 460226
rect 528390 460126 528514 460226
rect 528614 460126 530760 460226
rect 527580 460002 530760 460126
rect 527580 459902 527618 460002
rect 527718 459902 527842 460002
rect 527942 459902 528066 460002
rect 528166 459902 528290 460002
rect 528390 459902 528514 460002
rect 528614 459902 530760 460002
rect 527580 459778 530760 459902
rect 527580 459678 527618 459778
rect 527718 459678 527842 459778
rect 527942 459678 528066 459778
rect 528166 459678 528290 459778
rect 528390 459678 528514 459778
rect 528614 459678 530760 459778
rect 527580 459554 530760 459678
rect 527580 459454 527618 459554
rect 527718 459454 527842 459554
rect 527942 459454 528066 459554
rect 528166 459454 528290 459554
rect 528390 459454 528514 459554
rect 528614 459454 530760 459554
rect 527580 459330 530760 459454
rect 527580 459230 527618 459330
rect 527718 459230 527842 459330
rect 527942 459230 528066 459330
rect 528166 459230 528290 459330
rect 528390 459230 528514 459330
rect 528614 459230 530760 459330
rect 527580 459106 530760 459230
rect 527580 459006 527618 459106
rect 527718 459006 527842 459106
rect 527942 459006 528066 459106
rect 528166 459006 528290 459106
rect 528390 459006 528514 459106
rect 528614 459006 530760 459106
rect 527580 458882 530760 459006
rect 527580 458782 527618 458882
rect 527718 458782 527842 458882
rect 527942 458782 528066 458882
rect 528166 458782 528290 458882
rect 528390 458782 528514 458882
rect 528614 458782 530760 458882
rect 527580 458658 530760 458782
rect 527580 458558 527618 458658
rect 527718 458558 527842 458658
rect 527942 458558 528066 458658
rect 528166 458558 528290 458658
rect 528390 458558 528514 458658
rect 528614 458558 530760 458658
rect 527580 458434 530760 458558
rect 527580 458334 527618 458434
rect 527718 458334 527842 458434
rect 527942 458334 528066 458434
rect 528166 458334 528290 458434
rect 528390 458334 528514 458434
rect 528614 458334 530760 458434
rect 527580 458210 530760 458334
rect 527580 458110 527618 458210
rect 527718 458110 527842 458210
rect 527942 458110 528066 458210
rect 528166 458110 528290 458210
rect 528390 458110 528514 458210
rect 528614 458110 530760 458210
rect 527580 457986 530760 458110
rect 527580 457886 527618 457986
rect 527718 457886 527842 457986
rect 527942 457886 528066 457986
rect 528166 457886 528290 457986
rect 528390 457886 528514 457986
rect 528614 457886 530760 457986
rect 527580 457762 530760 457886
rect 527580 457662 527618 457762
rect 527718 457662 527842 457762
rect 527942 457662 528066 457762
rect 528166 457662 528290 457762
rect 528390 457662 528514 457762
rect 528614 457662 530760 457762
rect 527580 457538 530760 457662
rect 527580 457438 527618 457538
rect 527718 457438 527842 457538
rect 527942 457438 528066 457538
rect 528166 457438 528290 457538
rect 528390 457438 528514 457538
rect 528614 457452 530760 457538
rect 536504 457452 537320 462236
rect 528614 457438 537320 457452
rect 527580 457314 537320 457438
rect 527580 457214 527618 457314
rect 527718 457214 527842 457314
rect 527942 457214 528066 457314
rect 528166 457214 528290 457314
rect 528390 457214 528514 457314
rect 528614 457214 537320 457314
rect 527580 457176 537320 457214
rect 583520 455628 584800 455740
rect 562380 455440 567480 455520
rect 562380 455360 562480 455440
rect 562560 455360 562640 455440
rect 562720 455360 562800 455440
rect 562880 455360 562960 455440
rect 563040 455360 563120 455440
rect 563200 455360 563280 455440
rect 563360 455360 563440 455440
rect 563520 455360 563600 455440
rect 563680 455360 563760 455440
rect 563840 455360 563920 455440
rect 564000 455360 564080 455440
rect 564160 455360 564240 455440
rect 564320 455360 564400 455440
rect 564480 455360 564560 455440
rect 564640 455360 564720 455440
rect 564800 455360 564880 455440
rect 564960 455360 565040 455440
rect 565120 455360 565200 455440
rect 565280 455360 565360 455440
rect 565440 455360 565520 455440
rect 565600 455360 565680 455440
rect 565760 455360 565840 455440
rect 565920 455360 566000 455440
rect 566080 455360 566160 455440
rect 566240 455360 566320 455440
rect 566400 455360 566480 455440
rect 566560 455360 566640 455440
rect 566720 455360 566800 455440
rect 566880 455360 566960 455440
rect 567040 455360 567120 455440
rect 567200 455360 567280 455440
rect 567360 455360 567480 455440
rect 562380 455280 567480 455360
rect 562380 455200 562480 455280
rect 562560 455200 562640 455280
rect 562720 455200 562800 455280
rect 562880 455200 562960 455280
rect 563040 455200 563120 455280
rect 563200 455200 563280 455280
rect 563360 455200 563440 455280
rect 563520 455200 563600 455280
rect 563680 455200 563760 455280
rect 563840 455200 563920 455280
rect 564000 455200 564080 455280
rect 564160 455200 564240 455280
rect 564320 455200 564400 455280
rect 564480 455200 564560 455280
rect 564640 455200 564720 455280
rect 564800 455200 564880 455280
rect 564960 455200 565040 455280
rect 565120 455200 565200 455280
rect 565280 455200 565360 455280
rect 565440 455200 565520 455280
rect 565600 455200 565680 455280
rect 565760 455200 565840 455280
rect 565920 455200 566000 455280
rect 566080 455200 566160 455280
rect 566240 455200 566320 455280
rect 566400 455200 566480 455280
rect 566560 455200 566640 455280
rect 566720 455200 566800 455280
rect 566880 455200 566960 455280
rect 567040 455200 567120 455280
rect 567200 455200 567280 455280
rect 567360 455200 567480 455280
rect 562380 455160 567480 455200
rect 572540 455440 577640 455520
rect 572540 455360 572640 455440
rect 572720 455360 572800 455440
rect 572880 455360 572960 455440
rect 573040 455360 573120 455440
rect 573200 455360 573280 455440
rect 573360 455360 573440 455440
rect 573520 455360 573600 455440
rect 573680 455360 573760 455440
rect 573840 455360 573920 455440
rect 574000 455360 574080 455440
rect 574160 455360 574240 455440
rect 574320 455360 574400 455440
rect 574480 455360 574560 455440
rect 574640 455360 574720 455440
rect 574800 455360 574880 455440
rect 574960 455360 575040 455440
rect 575120 455360 575200 455440
rect 575280 455360 575360 455440
rect 575440 455360 575520 455440
rect 575600 455360 575680 455440
rect 575760 455360 575840 455440
rect 575920 455360 576000 455440
rect 576080 455360 576160 455440
rect 576240 455360 576320 455440
rect 576400 455360 576480 455440
rect 576560 455360 576640 455440
rect 576720 455360 576800 455440
rect 576880 455360 576960 455440
rect 577040 455360 577120 455440
rect 577200 455360 577280 455440
rect 577360 455360 577440 455440
rect 577520 455360 577640 455440
rect 572540 455280 577640 455360
rect 572540 455200 572640 455280
rect 572720 455200 572800 455280
rect 572880 455200 572960 455280
rect 573040 455200 573120 455280
rect 573200 455200 573280 455280
rect 573360 455200 573440 455280
rect 573520 455200 573600 455280
rect 573680 455200 573760 455280
rect 573840 455200 573920 455280
rect 574000 455200 574080 455280
rect 574160 455200 574240 455280
rect 574320 455200 574400 455280
rect 574480 455200 574560 455280
rect 574640 455200 574720 455280
rect 574800 455200 574880 455280
rect 574960 455200 575040 455280
rect 575120 455200 575200 455280
rect 575280 455200 575360 455280
rect 575440 455200 575520 455280
rect 575600 455200 575680 455280
rect 575760 455200 575840 455280
rect 575920 455200 576000 455280
rect 576080 455200 576160 455280
rect 576240 455200 576320 455280
rect 576400 455200 576480 455280
rect 576560 455200 576640 455280
rect 576720 455200 576800 455280
rect 576880 455200 576960 455280
rect 577040 455200 577120 455280
rect 577200 455200 577280 455280
rect 577360 455200 577440 455280
rect 577520 455200 577640 455280
rect 572540 455160 577640 455200
rect 583520 454446 584800 454558
rect 536120 454156 542702 454162
rect 512223 439877 513217 439882
rect 513520 453934 582788 454156
rect 513520 453919 572332 453934
rect 513520 453859 562222 453919
rect 562282 453859 562342 453919
rect 562402 453859 562462 453919
rect 562522 453859 562582 453919
rect 562642 453859 562702 453919
rect 562762 453859 562822 453919
rect 562882 453859 562942 453919
rect 563002 453859 563062 453919
rect 563122 453859 563182 453919
rect 563242 453859 563302 453919
rect 563362 453859 563422 453919
rect 563482 453859 563542 453919
rect 563602 453859 563662 453919
rect 563722 453859 563782 453919
rect 563842 453859 563902 453919
rect 563962 453859 564022 453919
rect 564082 453859 564142 453919
rect 564202 453859 564262 453919
rect 564322 453859 564382 453919
rect 564442 453859 564502 453919
rect 564562 453859 564622 453919
rect 564682 453859 564742 453919
rect 564802 453859 564862 453919
rect 564922 453859 564982 453919
rect 565042 453859 565102 453919
rect 565162 453859 565222 453919
rect 565282 453859 565342 453919
rect 565402 453859 565462 453919
rect 565522 453859 565582 453919
rect 565642 453859 565702 453919
rect 565762 453859 565822 453919
rect 565882 453859 565942 453919
rect 566002 453859 566062 453919
rect 566122 453859 566182 453919
rect 566242 453859 566302 453919
rect 566362 453859 566422 453919
rect 566482 453859 566542 453919
rect 566602 453859 566662 453919
rect 566722 453859 566782 453919
rect 566842 453859 566902 453919
rect 566962 453859 567022 453919
rect 567082 453859 567142 453919
rect 567202 453859 567262 453919
rect 567322 453859 567382 453919
rect 567442 453859 567502 453919
rect 567562 453874 572332 453919
rect 572392 453874 572452 453934
rect 572512 453874 572572 453934
rect 572632 453874 572692 453934
rect 572752 453874 572812 453934
rect 572872 453874 572932 453934
rect 572992 453874 573052 453934
rect 573112 453874 573172 453934
rect 573232 453874 573292 453934
rect 573352 453874 573412 453934
rect 573472 453874 573532 453934
rect 573592 453874 573652 453934
rect 573712 453874 573772 453934
rect 573832 453874 573892 453934
rect 573952 453874 574012 453934
rect 574072 453874 574132 453934
rect 574192 453874 574252 453934
rect 574312 453874 574372 453934
rect 574432 453874 574492 453934
rect 574552 453874 574612 453934
rect 574672 453874 574732 453934
rect 574792 453874 574852 453934
rect 574912 453874 574972 453934
rect 575032 453874 575092 453934
rect 575152 453874 575212 453934
rect 575272 453874 575332 453934
rect 575392 453874 575452 453934
rect 575512 453874 575572 453934
rect 575632 453874 575692 453934
rect 575752 453874 575812 453934
rect 575872 453874 575932 453934
rect 575992 453874 576052 453934
rect 576112 453874 576172 453934
rect 576232 453874 576292 453934
rect 576352 453874 576412 453934
rect 576472 453874 576532 453934
rect 576592 453874 576652 453934
rect 576712 453874 576772 453934
rect 576832 453874 576892 453934
rect 576952 453874 577012 453934
rect 577072 453874 577132 453934
rect 577192 453874 577252 453934
rect 577312 453874 577372 453934
rect 577432 453874 577492 453934
rect 577552 453874 577612 453934
rect 577672 453874 582788 453934
rect 567562 453859 582788 453874
rect 513520 453814 582788 453859
rect 513520 453799 572332 453814
rect 513520 453756 562222 453799
rect 513520 453556 513720 453756
rect 513920 453556 514154 453756
rect 514354 453556 514588 453756
rect 514788 453739 562222 453756
rect 562282 453739 562342 453799
rect 562402 453739 562462 453799
rect 562522 453739 562582 453799
rect 562642 453739 562702 453799
rect 562762 453739 562822 453799
rect 562882 453739 562942 453799
rect 563002 453739 563062 453799
rect 563122 453739 563182 453799
rect 563242 453739 563302 453799
rect 563362 453739 563422 453799
rect 563482 453739 563542 453799
rect 563602 453739 563662 453799
rect 563722 453739 563782 453799
rect 563842 453739 563902 453799
rect 563962 453739 564022 453799
rect 564082 453739 564142 453799
rect 564202 453739 564262 453799
rect 564322 453739 564382 453799
rect 564442 453739 564502 453799
rect 564562 453739 564622 453799
rect 564682 453739 564742 453799
rect 564802 453739 564862 453799
rect 564922 453739 564982 453799
rect 565042 453739 565102 453799
rect 565162 453739 565222 453799
rect 565282 453739 565342 453799
rect 565402 453739 565462 453799
rect 565522 453739 565582 453799
rect 565642 453739 565702 453799
rect 565762 453739 565822 453799
rect 565882 453739 565942 453799
rect 566002 453739 566062 453799
rect 566122 453739 566182 453799
rect 566242 453739 566302 453799
rect 566362 453739 566422 453799
rect 566482 453739 566542 453799
rect 566602 453739 566662 453799
rect 566722 453739 566782 453799
rect 566842 453739 566902 453799
rect 566962 453739 567022 453799
rect 567082 453739 567142 453799
rect 567202 453739 567262 453799
rect 567322 453739 567382 453799
rect 567442 453739 567502 453799
rect 567562 453754 572332 453799
rect 572392 453754 572452 453814
rect 572512 453754 572572 453814
rect 572632 453754 572692 453814
rect 572752 453754 572812 453814
rect 572872 453754 572932 453814
rect 572992 453754 573052 453814
rect 573112 453754 573172 453814
rect 573232 453754 573292 453814
rect 573352 453754 573412 453814
rect 573472 453754 573532 453814
rect 573592 453754 573652 453814
rect 573712 453754 573772 453814
rect 573832 453754 573892 453814
rect 573952 453754 574012 453814
rect 574072 453754 574132 453814
rect 574192 453754 574252 453814
rect 574312 453754 574372 453814
rect 574432 453754 574492 453814
rect 574552 453754 574612 453814
rect 574672 453754 574732 453814
rect 574792 453754 574852 453814
rect 574912 453754 574972 453814
rect 575032 453754 575092 453814
rect 575152 453754 575212 453814
rect 575272 453754 575332 453814
rect 575392 453754 575452 453814
rect 575512 453754 575572 453814
rect 575632 453754 575692 453814
rect 575752 453754 575812 453814
rect 575872 453754 575932 453814
rect 575992 453754 576052 453814
rect 576112 453754 576172 453814
rect 576232 453754 576292 453814
rect 576352 453754 576412 453814
rect 576472 453754 576532 453814
rect 576592 453754 576652 453814
rect 576712 453754 576772 453814
rect 576832 453754 576892 453814
rect 576952 453754 577012 453814
rect 577072 453754 577132 453814
rect 577192 453754 577252 453814
rect 577312 453754 577372 453814
rect 577432 453754 577492 453814
rect 577552 453754 577612 453814
rect 577672 453754 582788 453814
rect 567562 453739 582788 453754
rect 514788 453556 582788 453739
rect 513520 453322 582788 453556
rect 513520 453122 513720 453322
rect 513920 453122 514154 453322
rect 514354 453122 514588 453322
rect 514788 453122 582788 453322
rect 583520 453264 584800 453376
rect 513520 452888 582788 453122
rect 513520 452688 513720 452888
rect 513920 452688 514154 452888
rect 514354 452688 514588 452888
rect 514788 452688 582788 452888
rect 513520 452454 582788 452688
rect 513520 452254 513720 452454
rect 513920 452254 514154 452454
rect 514354 452254 514588 452454
rect 514788 452254 582788 452454
rect 513520 452020 582788 452254
rect 583520 452082 584800 452194
rect 513520 451820 513720 452020
rect 513920 451820 514154 452020
rect 514354 451820 514588 452020
rect 514788 451820 582788 452020
rect 513520 451586 582788 451820
rect 513520 451386 513720 451586
rect 513920 451386 514154 451586
rect 514354 451386 514588 451586
rect 514788 451386 582788 451586
rect 513520 451152 582788 451386
rect 513520 450952 513720 451152
rect 513920 450952 514154 451152
rect 514354 450952 514588 451152
rect 514788 450952 582788 451152
rect 513520 450718 582788 450952
rect 583520 450900 584800 451012
rect 513520 450518 513720 450718
rect 513920 450518 514154 450718
rect 514354 450518 514588 450718
rect 514788 450518 582788 450718
rect 513520 450284 582788 450518
rect 513520 450084 513720 450284
rect 513920 450084 514154 450284
rect 514354 450084 514588 450284
rect 514788 450084 582788 450284
rect 513520 449850 582788 450084
rect 513520 449650 513720 449850
rect 513920 449650 514154 449850
rect 514354 449650 514588 449850
rect 514788 449830 582788 449850
rect 514788 449718 584800 449830
rect 514788 449650 582788 449718
rect 513520 449416 582788 449650
rect 513520 449216 513720 449416
rect 513920 449216 514154 449416
rect 514354 449216 514588 449416
rect 514788 449216 582788 449416
rect 513520 449016 582788 449216
rect 513520 448816 514588 449016
rect 514788 448816 582788 449016
rect 513520 448616 582788 448816
rect 513520 448416 514588 448616
rect 514788 448416 582788 448616
rect 513520 448216 582788 448416
rect 513520 448016 514588 448216
rect 514788 448016 582788 448216
rect 513520 447816 582788 448016
rect 513520 447616 514588 447816
rect 514788 447616 582788 447816
rect 513520 447416 582788 447616
rect 513520 447216 514588 447416
rect 514788 447216 582788 447416
rect 513520 447016 582788 447216
rect 513520 446816 514588 447016
rect 514788 446816 582788 447016
rect 513520 446616 582788 446816
rect 513520 446416 514588 446616
rect 514788 446416 582788 446616
rect 513520 446216 582788 446416
rect 513520 446016 514588 446216
rect 514788 446016 582788 446216
rect 513520 445816 582788 446016
rect 513520 445616 514588 445816
rect 514788 445616 582788 445816
rect 513520 444216 582788 445616
rect 513520 444016 514588 444216
rect 514788 444016 582788 444216
rect 513520 443816 582788 444016
rect 513520 443616 514588 443816
rect 514788 443616 582788 443816
rect 513520 443416 582788 443616
rect 513520 443216 514588 443416
rect 514788 443216 582788 443416
rect 513520 443016 582788 443216
rect 513520 442816 514588 443016
rect 514788 442816 582788 443016
rect 513520 442616 582788 442816
rect 513520 442416 514588 442616
rect 514788 442416 582788 442616
rect 513520 442216 582788 442416
rect 513520 442016 514588 442216
rect 514788 442016 582788 442216
rect 513520 441816 582788 442016
rect 513520 441616 514588 441816
rect 514788 441616 582788 441816
rect 513520 441416 582788 441616
rect 513520 441216 514588 441416
rect 514788 441216 582788 441416
rect 513520 441016 582788 441216
rect 513520 440816 514588 441016
rect 514788 440816 582788 441016
rect 513520 438756 582788 440816
rect 500384 437576 501460 437596
rect 527604 437576 528664 437580
rect 490640 437540 501460 437576
rect 490640 437440 500418 437540
rect 500518 437440 500642 437540
rect 500742 437440 500866 437540
rect 500966 437440 501090 437540
rect 501190 437440 501314 437540
rect 501414 437440 501460 437540
rect 490640 437316 501460 437440
rect 490640 437216 500418 437316
rect 500518 437216 500642 437316
rect 500742 437216 500866 437316
rect 500966 437216 501090 437316
rect 501190 437216 501314 437316
rect 501414 437216 501460 437316
rect 490640 437092 501460 437216
rect 490640 436992 500418 437092
rect 500518 436992 500642 437092
rect 500742 436992 500866 437092
rect 500966 436992 501090 437092
rect 501190 436992 501314 437092
rect 501414 436992 501460 437092
rect 490640 436868 501460 436992
rect 490640 436768 500418 436868
rect 500518 436768 500642 436868
rect 500742 436768 500866 436868
rect 500966 436768 501090 436868
rect 501190 436768 501314 436868
rect 501414 436768 501460 436868
rect 490640 436676 501460 436768
rect 490640 431892 491260 436676
rect 497004 436644 501460 436676
rect 497004 436544 500418 436644
rect 500518 436544 500642 436644
rect 500742 436544 500866 436644
rect 500966 436544 501090 436644
rect 501190 436544 501314 436644
rect 501414 436544 501460 436644
rect 497004 436420 501460 436544
rect 497004 436320 500418 436420
rect 500518 436320 500642 436420
rect 500742 436320 500866 436420
rect 500966 436320 501090 436420
rect 501190 436320 501314 436420
rect 501414 436320 501460 436420
rect 497004 436196 501460 436320
rect 497004 436096 500418 436196
rect 500518 436096 500642 436196
rect 500742 436096 500866 436196
rect 500966 436096 501090 436196
rect 501190 436096 501314 436196
rect 501414 436096 501460 436196
rect 497004 435972 501460 436096
rect 497004 435872 500418 435972
rect 500518 435872 500642 435972
rect 500742 435872 500866 435972
rect 500966 435872 501090 435972
rect 501190 435872 501314 435972
rect 501414 435872 501460 435972
rect 497004 435748 501460 435872
rect 497004 435648 500418 435748
rect 500518 435648 500642 435748
rect 500742 435648 500866 435748
rect 500966 435648 501090 435748
rect 501190 435648 501314 435748
rect 501414 435648 501460 435748
rect 497004 435524 501460 435648
rect 497004 435424 500418 435524
rect 500518 435424 500642 435524
rect 500742 435424 500866 435524
rect 500966 435424 501090 435524
rect 501190 435424 501314 435524
rect 501414 435424 501460 435524
rect 497004 435300 501460 435424
rect 497004 435200 500418 435300
rect 500518 435200 500642 435300
rect 500742 435200 500866 435300
rect 500966 435200 501090 435300
rect 501190 435200 501314 435300
rect 501414 435200 501460 435300
rect 497004 435076 501460 435200
rect 497004 434976 500418 435076
rect 500518 434976 500642 435076
rect 500742 434976 500866 435076
rect 500966 434976 501090 435076
rect 501190 434976 501314 435076
rect 501414 434976 501460 435076
rect 497004 434852 501460 434976
rect 497004 434752 500418 434852
rect 500518 434752 500642 434852
rect 500742 434752 500866 434852
rect 500966 434752 501090 434852
rect 501190 434752 501314 434852
rect 501414 434752 501460 434852
rect 497004 434628 501460 434752
rect 497004 434528 500418 434628
rect 500518 434528 500642 434628
rect 500742 434528 500866 434628
rect 500966 434528 501090 434628
rect 501190 434528 501314 434628
rect 501414 434528 501460 434628
rect 497004 434404 501460 434528
rect 497004 434304 500418 434404
rect 500518 434304 500642 434404
rect 500742 434304 500866 434404
rect 500966 434304 501090 434404
rect 501190 434304 501314 434404
rect 501414 434304 501460 434404
rect 497004 434180 501460 434304
rect 497004 434080 500418 434180
rect 500518 434080 500642 434180
rect 500742 434080 500866 434180
rect 500966 434080 501090 434180
rect 501190 434080 501314 434180
rect 501414 434080 501460 434180
rect 497004 433956 501460 434080
rect 497004 433856 500418 433956
rect 500518 433856 500642 433956
rect 500742 433856 500866 433956
rect 500966 433856 501090 433956
rect 501190 433856 501314 433956
rect 501414 433856 501460 433956
rect 497004 433732 501460 433856
rect 497004 433632 500418 433732
rect 500518 433632 500642 433732
rect 500742 433632 500866 433732
rect 500966 433632 501090 433732
rect 501190 433632 501314 433732
rect 501414 433632 501460 433732
rect 497004 433508 501460 433632
rect 497004 433408 500418 433508
rect 500518 433408 500642 433508
rect 500742 433408 500866 433508
rect 500966 433408 501090 433508
rect 501190 433408 501314 433508
rect 501414 433408 501460 433508
rect 497004 433284 501460 433408
rect 497004 433184 500418 433284
rect 500518 433184 500642 433284
rect 500742 433184 500866 433284
rect 500966 433184 501090 433284
rect 501190 433184 501314 433284
rect 501414 433184 501460 433284
rect 497004 433060 501460 433184
rect 497004 432960 500418 433060
rect 500518 432960 500642 433060
rect 500742 432960 500866 433060
rect 500966 432960 501090 433060
rect 501190 432960 501314 433060
rect 501414 432960 501460 433060
rect 497004 432836 501460 432960
rect 497004 432736 500418 432836
rect 500518 432736 500642 432836
rect 500742 432736 500866 432836
rect 500966 432736 501090 432836
rect 501190 432736 501314 432836
rect 501414 432736 501460 432836
rect 497004 432612 501460 432736
rect 497004 432512 500418 432612
rect 500518 432512 500642 432612
rect 500742 432512 500866 432612
rect 500966 432512 501090 432612
rect 501190 432512 501314 432612
rect 501414 432512 501460 432612
rect 497004 432388 501460 432512
rect 497004 432288 500418 432388
rect 500518 432288 500642 432388
rect 500742 432288 500866 432388
rect 500966 432288 501090 432388
rect 501190 432288 501314 432388
rect 501414 432288 501460 432388
rect 497004 432164 501460 432288
rect 497004 432064 500418 432164
rect 500518 432064 500642 432164
rect 500742 432064 500866 432164
rect 500966 432064 501090 432164
rect 501190 432064 501314 432164
rect 501414 432064 501460 432164
rect 497004 431940 501460 432064
rect 497004 431892 500418 431940
rect 490640 431840 500418 431892
rect 500518 431840 500642 431940
rect 500742 431840 500866 431940
rect 500966 431840 501090 431940
rect 501190 431840 501314 431940
rect 501414 431840 501460 431940
rect 490640 431716 501460 431840
rect 490640 431616 500418 431716
rect 500518 431616 500642 431716
rect 500742 431616 500866 431716
rect 500966 431616 501090 431716
rect 501190 431616 501314 431716
rect 501414 431616 501460 431716
rect 490640 431492 501460 431616
rect 490640 431392 500418 431492
rect 500518 431392 500642 431492
rect 500742 431392 500866 431492
rect 500966 431392 501090 431492
rect 501190 431392 501314 431492
rect 501414 431392 501460 431492
rect 490640 431268 501460 431392
rect 490640 431168 500418 431268
rect 500518 431168 500642 431268
rect 500742 431168 500866 431268
rect 500966 431168 501090 431268
rect 501190 431168 501314 431268
rect 501414 431168 501460 431268
rect 490640 431044 501460 431168
rect 527580 437540 537300 437576
rect 527580 437440 527638 437540
rect 527738 437440 527862 437540
rect 527962 437440 528086 437540
rect 528186 437440 528310 437540
rect 528410 437440 528534 437540
rect 528634 437440 537300 437540
rect 527580 437316 537300 437440
rect 527580 437216 527638 437316
rect 527738 437216 527862 437316
rect 527962 437216 528086 437316
rect 528186 437216 528310 437316
rect 528410 437216 528534 437316
rect 528634 437216 537300 437316
rect 527580 437092 537300 437216
rect 527580 436992 527638 437092
rect 527738 436992 527862 437092
rect 527962 436992 528086 437092
rect 528186 436992 528310 437092
rect 528410 436992 528534 437092
rect 528634 436992 537300 437092
rect 527580 436868 537300 436992
rect 527580 436768 527638 436868
rect 527738 436768 527862 436868
rect 527962 436768 528086 436868
rect 528186 436768 528310 436868
rect 528410 436768 528534 436868
rect 528634 436768 537300 436868
rect 527580 436676 537300 436768
rect 527580 436644 531080 436676
rect 527580 436544 527638 436644
rect 527738 436544 527862 436644
rect 527962 436544 528086 436644
rect 528186 436544 528310 436644
rect 528410 436544 528534 436644
rect 528634 436544 531080 436644
rect 527580 436420 531080 436544
rect 527580 436320 527638 436420
rect 527738 436320 527862 436420
rect 527962 436320 528086 436420
rect 528186 436320 528310 436420
rect 528410 436320 528534 436420
rect 528634 436320 531080 436420
rect 527580 436196 531080 436320
rect 527580 436096 527638 436196
rect 527738 436096 527862 436196
rect 527962 436096 528086 436196
rect 528186 436096 528310 436196
rect 528410 436096 528534 436196
rect 528634 436096 531080 436196
rect 527580 435972 531080 436096
rect 527580 435872 527638 435972
rect 527738 435872 527862 435972
rect 527962 435872 528086 435972
rect 528186 435872 528310 435972
rect 528410 435872 528534 435972
rect 528634 435872 531080 435972
rect 527580 435748 531080 435872
rect 527580 435648 527638 435748
rect 527738 435648 527862 435748
rect 527962 435648 528086 435748
rect 528186 435648 528310 435748
rect 528410 435648 528534 435748
rect 528634 435648 531080 435748
rect 527580 435524 531080 435648
rect 527580 435424 527638 435524
rect 527738 435424 527862 435524
rect 527962 435424 528086 435524
rect 528186 435424 528310 435524
rect 528410 435424 528534 435524
rect 528634 435424 531080 435524
rect 527580 435300 531080 435424
rect 527580 435200 527638 435300
rect 527738 435200 527862 435300
rect 527962 435200 528086 435300
rect 528186 435200 528310 435300
rect 528410 435200 528534 435300
rect 528634 435200 531080 435300
rect 527580 435076 531080 435200
rect 527580 434976 527638 435076
rect 527738 434976 527862 435076
rect 527962 434976 528086 435076
rect 528186 434976 528310 435076
rect 528410 434976 528534 435076
rect 528634 434976 531080 435076
rect 527580 434852 531080 434976
rect 527580 434752 527638 434852
rect 527738 434752 527862 434852
rect 527962 434752 528086 434852
rect 528186 434752 528310 434852
rect 528410 434752 528534 434852
rect 528634 434752 531080 434852
rect 527580 434628 531080 434752
rect 527580 434528 527638 434628
rect 527738 434528 527862 434628
rect 527962 434528 528086 434628
rect 528186 434528 528310 434628
rect 528410 434528 528534 434628
rect 528634 434528 531080 434628
rect 527580 434404 531080 434528
rect 527580 434304 527638 434404
rect 527738 434304 527862 434404
rect 527962 434304 528086 434404
rect 528186 434304 528310 434404
rect 528410 434304 528534 434404
rect 528634 434304 531080 434404
rect 527580 434180 531080 434304
rect 527580 434080 527638 434180
rect 527738 434080 527862 434180
rect 527962 434080 528086 434180
rect 528186 434080 528310 434180
rect 528410 434080 528534 434180
rect 528634 434080 531080 434180
rect 527580 433956 531080 434080
rect 527580 433856 527638 433956
rect 527738 433856 527862 433956
rect 527962 433856 528086 433956
rect 528186 433856 528310 433956
rect 528410 433856 528534 433956
rect 528634 433856 531080 433956
rect 527580 433732 531080 433856
rect 527580 433632 527638 433732
rect 527738 433632 527862 433732
rect 527962 433632 528086 433732
rect 528186 433632 528310 433732
rect 528410 433632 528534 433732
rect 528634 433632 531080 433732
rect 527580 433508 531080 433632
rect 527580 433408 527638 433508
rect 527738 433408 527862 433508
rect 527962 433408 528086 433508
rect 528186 433408 528310 433508
rect 528410 433408 528534 433508
rect 528634 433408 531080 433508
rect 527580 433284 531080 433408
rect 527580 433184 527638 433284
rect 527738 433184 527862 433284
rect 527962 433184 528086 433284
rect 528186 433184 528310 433284
rect 528410 433184 528534 433284
rect 528634 433184 531080 433284
rect 527580 433060 531080 433184
rect 527580 432960 527638 433060
rect 527738 432960 527862 433060
rect 527962 432960 528086 433060
rect 528186 432960 528310 433060
rect 528410 432960 528534 433060
rect 528634 432960 531080 433060
rect 527580 432836 531080 432960
rect 527580 432736 527638 432836
rect 527738 432736 527862 432836
rect 527962 432736 528086 432836
rect 528186 432736 528310 432836
rect 528410 432736 528534 432836
rect 528634 432736 531080 432836
rect 527580 432612 531080 432736
rect 527580 432512 527638 432612
rect 527738 432512 527862 432612
rect 527962 432512 528086 432612
rect 528186 432512 528310 432612
rect 528410 432512 528534 432612
rect 528634 432512 531080 432612
rect 527580 432388 531080 432512
rect 527580 432288 527638 432388
rect 527738 432288 527862 432388
rect 527962 432288 528086 432388
rect 528186 432288 528310 432388
rect 528410 432288 528534 432388
rect 528634 432288 531080 432388
rect 527580 432164 531080 432288
rect 527580 432064 527638 432164
rect 527738 432064 527862 432164
rect 527962 432064 528086 432164
rect 528186 432064 528310 432164
rect 528410 432064 528534 432164
rect 528634 432064 531080 432164
rect 527580 431940 531080 432064
rect 527580 431840 527638 431940
rect 527738 431840 527862 431940
rect 527962 431840 528086 431940
rect 528186 431840 528310 431940
rect 528410 431840 528534 431940
rect 528634 431892 531080 431940
rect 536824 431892 537300 436676
rect 528634 431840 537300 431892
rect 527580 431716 537300 431840
rect 527580 431616 527638 431716
rect 527738 431616 527862 431716
rect 527962 431616 528086 431716
rect 528186 431616 528310 431716
rect 528410 431616 528534 431716
rect 528634 431616 537300 431716
rect 527580 431492 537300 431616
rect 527580 431392 527638 431492
rect 527738 431392 527862 431492
rect 527962 431392 528086 431492
rect 528186 431392 528310 431492
rect 528410 431392 528534 431492
rect 528634 431392 537300 431492
rect 527580 431268 537300 431392
rect 527580 431168 527638 431268
rect 527738 431168 527862 431268
rect 527962 431168 528086 431268
rect 528186 431168 528310 431268
rect 528410 431168 528534 431268
rect 528634 431168 537300 431268
rect 490640 430944 500418 431044
rect 500518 430944 500642 431044
rect 500742 430944 500866 431044
rect 500966 430944 501090 431044
rect 501190 430944 501314 431044
rect 501414 430944 501460 431044
rect 490640 430756 501460 430944
rect 503864 431056 510520 431156
rect 503864 431026 510526 431056
rect 503864 430926 503920 431026
rect 504020 430926 504144 431026
rect 504244 430926 504368 431026
rect 504468 430926 504592 431026
rect 504692 430926 504816 431026
rect 504916 430926 505040 431026
rect 505140 430926 505264 431026
rect 505364 430926 505488 431026
rect 505588 430926 505712 431026
rect 505812 430926 505936 431026
rect 506036 430926 506160 431026
rect 506260 430926 506384 431026
rect 506484 430926 506608 431026
rect 506708 430926 506832 431026
rect 506932 430926 507056 431026
rect 507156 430926 507280 431026
rect 507380 430926 507504 431026
rect 507604 430926 507728 431026
rect 507828 430926 507952 431026
rect 508052 430926 508176 431026
rect 508276 430926 508400 431026
rect 508500 430926 508624 431026
rect 508724 430926 508848 431026
rect 508948 430926 509072 431026
rect 509172 430926 509296 431026
rect 509396 430926 509520 431026
rect 509620 430926 509744 431026
rect 509844 430926 509968 431026
rect 510068 430926 510192 431026
rect 510292 430926 510416 431026
rect 510516 430926 510526 431026
rect 503864 430802 510526 430926
rect 503864 430702 503920 430802
rect 504020 430702 504144 430802
rect 504244 430702 504368 430802
rect 504468 430702 504592 430802
rect 504692 430702 504816 430802
rect 504916 430702 505040 430802
rect 505140 430702 505264 430802
rect 505364 430702 505488 430802
rect 505588 430702 505712 430802
rect 505812 430702 505936 430802
rect 506036 430702 506160 430802
rect 506260 430702 506384 430802
rect 506484 430702 506608 430802
rect 506708 430702 506832 430802
rect 506932 430702 507056 430802
rect 507156 430702 507280 430802
rect 507380 430702 507504 430802
rect 507604 430702 507728 430802
rect 507828 430702 507952 430802
rect 508052 430702 508176 430802
rect 508276 430702 508400 430802
rect 508500 430702 508624 430802
rect 508724 430702 508848 430802
rect 508948 430702 509072 430802
rect 509172 430702 509296 430802
rect 509396 430702 509520 430802
rect 509620 430702 509744 430802
rect 509844 430702 509968 430802
rect 510068 430702 510192 430802
rect 510292 430702 510416 430802
rect 510516 430702 510526 430802
rect 503864 430578 510526 430702
rect 503864 430478 503920 430578
rect 504020 430478 504144 430578
rect 504244 430478 504368 430578
rect 504468 430478 504592 430578
rect 504692 430478 504816 430578
rect 504916 430478 505040 430578
rect 505140 430478 505264 430578
rect 505364 430478 505488 430578
rect 505588 430478 505712 430578
rect 505812 430478 505936 430578
rect 506036 430478 506160 430578
rect 506260 430478 506384 430578
rect 506484 430478 506608 430578
rect 506708 430478 506832 430578
rect 506932 430478 507056 430578
rect 507156 430478 507280 430578
rect 507380 430478 507504 430578
rect 507604 430478 507728 430578
rect 507828 430478 507952 430578
rect 508052 430478 508176 430578
rect 508276 430478 508400 430578
rect 508500 430478 508624 430578
rect 508724 430478 508848 430578
rect 508948 430478 509072 430578
rect 509172 430478 509296 430578
rect 509396 430478 509520 430578
rect 509620 430478 509744 430578
rect 509844 430478 509968 430578
rect 510068 430478 510192 430578
rect 510292 430478 510416 430578
rect 510516 430478 510526 430578
rect 503864 430354 510526 430478
rect 503864 430254 503920 430354
rect 504020 430254 504144 430354
rect 504244 430254 504368 430354
rect 504468 430254 504592 430354
rect 504692 430254 504816 430354
rect 504916 430254 505040 430354
rect 505140 430254 505264 430354
rect 505364 430254 505488 430354
rect 505588 430254 505712 430354
rect 505812 430254 505936 430354
rect 506036 430254 506160 430354
rect 506260 430254 506384 430354
rect 506484 430254 506608 430354
rect 506708 430254 506832 430354
rect 506932 430254 507056 430354
rect 507156 430254 507280 430354
rect 507380 430254 507504 430354
rect 507604 430254 507728 430354
rect 507828 430254 507952 430354
rect 508052 430254 508176 430354
rect 508276 430254 508400 430354
rect 508500 430254 508624 430354
rect 508724 430254 508848 430354
rect 508948 430254 509072 430354
rect 509172 430254 509296 430354
rect 509396 430254 509520 430354
rect 509620 430254 509744 430354
rect 509844 430254 509968 430354
rect 510068 430254 510192 430354
rect 510292 430254 510416 430354
rect 510516 430254 510526 430354
rect 503864 430130 510526 430254
rect 503864 430030 503920 430130
rect 504020 430030 504144 430130
rect 504244 430030 504368 430130
rect 504468 430030 504592 430130
rect 504692 430030 504816 430130
rect 504916 430030 505040 430130
rect 505140 430030 505264 430130
rect 505364 430030 505488 430130
rect 505588 430030 505712 430130
rect 505812 430030 505936 430130
rect 506036 430030 506160 430130
rect 506260 430030 506384 430130
rect 506484 430030 506608 430130
rect 506708 430030 506832 430130
rect 506932 430030 507056 430130
rect 507156 430030 507280 430130
rect 507380 430030 507504 430130
rect 507604 430030 507728 430130
rect 507828 430030 507952 430130
rect 508052 430030 508176 430130
rect 508276 430030 508400 430130
rect 508500 430030 508624 430130
rect 508724 430030 508848 430130
rect 508948 430030 509072 430130
rect 509172 430030 509296 430130
rect 509396 430030 509520 430130
rect 509620 430030 509744 430130
rect 509844 430030 509968 430130
rect 510068 430030 510192 430130
rect 510292 430030 510416 430130
rect 510516 430030 510526 430130
rect 503864 429970 510526 430030
rect 517280 431026 523940 431056
rect 517280 430926 517320 431026
rect 517420 430926 517544 431026
rect 517644 430926 517768 431026
rect 517868 430926 517992 431026
rect 518092 430926 518216 431026
rect 518316 430926 518440 431026
rect 518540 430926 518664 431026
rect 518764 430926 518888 431026
rect 518988 430926 519112 431026
rect 519212 430926 519336 431026
rect 519436 430926 519560 431026
rect 519660 430926 519784 431026
rect 519884 430926 520008 431026
rect 520108 430926 520232 431026
rect 520332 430926 520456 431026
rect 520556 430926 520680 431026
rect 520780 430926 520904 431026
rect 521004 430926 521128 431026
rect 521228 430926 521352 431026
rect 521452 430926 521576 431026
rect 521676 430926 521800 431026
rect 521900 430926 522024 431026
rect 522124 430926 522248 431026
rect 522348 430926 522472 431026
rect 522572 430926 522696 431026
rect 522796 430926 522920 431026
rect 523020 430926 523144 431026
rect 523244 430926 523368 431026
rect 523468 430926 523592 431026
rect 523692 430926 523816 431026
rect 523916 430926 523940 431026
rect 517280 430802 523940 430926
rect 517280 430702 517320 430802
rect 517420 430702 517544 430802
rect 517644 430702 517768 430802
rect 517868 430702 517992 430802
rect 518092 430702 518216 430802
rect 518316 430702 518440 430802
rect 518540 430702 518664 430802
rect 518764 430702 518888 430802
rect 518988 430702 519112 430802
rect 519212 430702 519336 430802
rect 519436 430702 519560 430802
rect 519660 430702 519784 430802
rect 519884 430702 520008 430802
rect 520108 430702 520232 430802
rect 520332 430702 520456 430802
rect 520556 430702 520680 430802
rect 520780 430702 520904 430802
rect 521004 430702 521128 430802
rect 521228 430702 521352 430802
rect 521452 430702 521576 430802
rect 521676 430702 521800 430802
rect 521900 430702 522024 430802
rect 522124 430702 522248 430802
rect 522348 430702 522472 430802
rect 522572 430702 522696 430802
rect 522796 430702 522920 430802
rect 523020 430702 523144 430802
rect 523244 430702 523368 430802
rect 523468 430702 523592 430802
rect 523692 430702 523816 430802
rect 523916 430702 523940 430802
rect 527580 431044 537300 431168
rect 527580 430944 527638 431044
rect 527738 430944 527862 431044
rect 527962 430944 528086 431044
rect 528186 430944 528310 431044
rect 528410 430944 528534 431044
rect 528634 430944 537300 431044
rect 527580 430756 537300 430944
rect 517280 430578 523940 430702
rect 517280 430478 517320 430578
rect 517420 430478 517544 430578
rect 517644 430478 517768 430578
rect 517868 430478 517992 430578
rect 518092 430478 518216 430578
rect 518316 430478 518440 430578
rect 518540 430478 518664 430578
rect 518764 430478 518888 430578
rect 518988 430478 519112 430578
rect 519212 430478 519336 430578
rect 519436 430478 519560 430578
rect 519660 430478 519784 430578
rect 519884 430478 520008 430578
rect 520108 430478 520232 430578
rect 520332 430478 520456 430578
rect 520556 430478 520680 430578
rect 520780 430478 520904 430578
rect 521004 430478 521128 430578
rect 521228 430478 521352 430578
rect 521452 430478 521576 430578
rect 521676 430478 521800 430578
rect 521900 430478 522024 430578
rect 522124 430478 522248 430578
rect 522348 430478 522472 430578
rect 522572 430478 522696 430578
rect 522796 430478 522920 430578
rect 523020 430478 523144 430578
rect 523244 430478 523368 430578
rect 523468 430478 523592 430578
rect 523692 430478 523816 430578
rect 523916 430478 523940 430578
rect 517280 430354 523940 430478
rect 517280 430254 517320 430354
rect 517420 430254 517544 430354
rect 517644 430254 517768 430354
rect 517868 430254 517992 430354
rect 518092 430254 518216 430354
rect 518316 430254 518440 430354
rect 518540 430254 518664 430354
rect 518764 430254 518888 430354
rect 518988 430254 519112 430354
rect 519212 430254 519336 430354
rect 519436 430254 519560 430354
rect 519660 430254 519784 430354
rect 519884 430254 520008 430354
rect 520108 430254 520232 430354
rect 520332 430254 520456 430354
rect 520556 430254 520680 430354
rect 520780 430254 520904 430354
rect 521004 430254 521128 430354
rect 521228 430254 521352 430354
rect 521452 430254 521576 430354
rect 521676 430254 521800 430354
rect 521900 430254 522024 430354
rect 522124 430254 522248 430354
rect 522348 430254 522472 430354
rect 522572 430254 522696 430354
rect 522796 430254 522920 430354
rect 523020 430254 523144 430354
rect 523244 430254 523368 430354
rect 523468 430254 523592 430354
rect 523692 430254 523816 430354
rect 523916 430254 523940 430354
rect 517280 430130 523940 430254
rect 517280 430030 517320 430130
rect 517420 430030 517544 430130
rect 517644 430030 517768 430130
rect 517868 430030 517992 430130
rect 518092 430030 518216 430130
rect 518316 430030 518440 430130
rect 518540 430030 518664 430130
rect 518764 430030 518888 430130
rect 518988 430030 519112 430130
rect 519212 430030 519336 430130
rect 519436 430030 519560 430130
rect 519660 430030 519784 430130
rect 519884 430030 520008 430130
rect 520108 430030 520232 430130
rect 520332 430030 520456 430130
rect 520556 430030 520680 430130
rect 520780 430030 520904 430130
rect 521004 430030 521128 430130
rect 521228 430030 521352 430130
rect 521452 430030 521576 430130
rect 521676 430030 521800 430130
rect 521900 430030 522024 430130
rect 522124 430030 522248 430130
rect 522348 430030 522472 430130
rect 522572 430030 522696 430130
rect 522796 430030 522920 430130
rect 523020 430030 523144 430130
rect 523244 430030 523368 430130
rect 523468 430030 523592 430130
rect 523692 430030 523816 430130
rect 523916 430030 523940 430130
rect 517280 429996 523940 430030
rect 490482 426452 578882 426928
rect 490482 426216 572772 426452
rect 573008 426216 573244 426452
rect 573480 426216 573716 426452
rect 573952 426216 574188 426452
rect 574424 426216 574660 426452
rect 574896 426216 575132 426452
rect 575368 426216 575604 426452
rect 575840 426216 576076 426452
rect 576312 426216 576548 426452
rect 576784 426216 577020 426452
rect 577256 426216 578882 426452
rect 490482 426000 578882 426216
rect -800 425086 480 425198
rect -800 423904 480 424016
rect -800 422722 480 422834
rect -800 421540 480 421652
rect 490482 421216 491138 426000
rect 496882 421216 504338 426000
rect 510082 421216 517738 426000
rect 523482 421216 531138 426000
rect 536882 425980 578882 426000
rect 536882 425744 572772 425980
rect 573008 425744 573244 425980
rect 573480 425744 573716 425980
rect 573952 425744 574188 425980
rect 574424 425744 574660 425980
rect 574896 425744 575132 425980
rect 575368 425744 575604 425980
rect 575840 425744 576076 425980
rect 576312 425744 576548 425980
rect 576784 425744 577020 425980
rect 577256 425744 578882 425980
rect 536882 425508 578882 425744
rect 536882 425272 572772 425508
rect 573008 425272 573244 425508
rect 573480 425272 573716 425508
rect 573952 425272 574188 425508
rect 574424 425272 574660 425508
rect 574896 425272 575132 425508
rect 575368 425272 575604 425508
rect 575840 425272 576076 425508
rect 576312 425272 576548 425508
rect 576784 425272 577020 425508
rect 577256 425272 578882 425508
rect 536882 425036 578882 425272
rect 536882 424800 572772 425036
rect 573008 424800 573244 425036
rect 573480 424800 573716 425036
rect 573952 424800 574188 425036
rect 574424 424800 574660 425036
rect 574896 424800 575132 425036
rect 575368 424800 575604 425036
rect 575840 424800 576076 425036
rect 576312 424800 576548 425036
rect 576784 424800 577020 425036
rect 577256 424800 578882 425036
rect 536882 424564 578882 424800
rect 536882 424328 572772 424564
rect 573008 424328 573244 424564
rect 573480 424328 573716 424564
rect 573952 424328 574188 424564
rect 574424 424328 574660 424564
rect 574896 424328 575132 424564
rect 575368 424328 575604 424564
rect 575840 424328 576076 424564
rect 576312 424328 576548 424564
rect 576784 424328 577020 424564
rect 577256 424328 578882 424564
rect 536882 424092 578882 424328
rect 536882 423856 572772 424092
rect 573008 423856 573244 424092
rect 573480 423856 573716 424092
rect 573952 423856 574188 424092
rect 574424 423856 574660 424092
rect 574896 423856 575132 424092
rect 575368 423856 575604 424092
rect 575840 423856 576076 424092
rect 576312 423856 576548 424092
rect 576784 423856 577020 424092
rect 577256 423856 578882 424092
rect 536882 423620 578882 423856
rect 536882 423384 572772 423620
rect 573008 423384 573244 423620
rect 573480 423384 573716 423620
rect 573952 423384 574188 423620
rect 574424 423384 574660 423620
rect 574896 423384 575132 423620
rect 575368 423384 575604 423620
rect 575840 423384 576076 423620
rect 576312 423384 576548 423620
rect 576784 423384 577020 423620
rect 577256 423384 578882 423620
rect 536882 423148 578882 423384
rect 536882 422912 572772 423148
rect 573008 422912 573244 423148
rect 573480 422912 573716 423148
rect 573952 422912 574188 423148
rect 574424 422912 574660 423148
rect 574896 422912 575132 423148
rect 575368 422912 575604 423148
rect 575840 422912 576076 423148
rect 576312 422912 576548 423148
rect 576784 422912 577020 423148
rect 577256 422912 578882 423148
rect 536882 422676 578882 422912
rect 536882 422440 572772 422676
rect 573008 422440 573244 422676
rect 573480 422440 573716 422676
rect 573952 422440 574188 422676
rect 574424 422440 574660 422676
rect 574896 422440 575132 422676
rect 575368 422440 575604 422676
rect 575840 422440 576076 422676
rect 576312 422440 576548 422676
rect 576784 422440 577020 422676
rect 577256 422440 578882 422676
rect 536882 422204 578882 422440
rect 536882 421968 572772 422204
rect 573008 421968 573244 422204
rect 573480 421968 573716 422204
rect 573952 421968 574188 422204
rect 574424 421968 574660 422204
rect 574896 421968 575132 422204
rect 575368 421968 575604 422204
rect 575840 421968 576076 422204
rect 576312 421968 576548 422204
rect 576784 421968 577020 422204
rect 577256 421968 578882 422204
rect 536882 421732 578882 421968
rect 536882 421496 572772 421732
rect 573008 421496 573244 421732
rect 573480 421496 573716 421732
rect 573952 421496 574188 421732
rect 574424 421496 574660 421732
rect 574896 421496 575132 421732
rect 575368 421496 575604 421732
rect 575840 421496 576076 421732
rect 576312 421496 576548 421732
rect 576784 421496 577020 421732
rect 577256 421496 578882 421732
rect 536882 421260 578882 421496
rect 536882 421216 572772 421260
rect 490482 421024 572772 421216
rect 573008 421024 573244 421260
rect 573480 421024 573716 421260
rect 573952 421024 574188 421260
rect 574424 421024 574660 421260
rect 574896 421024 575132 421260
rect 575368 421024 575604 421260
rect 575840 421024 576076 421260
rect 576312 421024 576548 421260
rect 576784 421024 577020 421260
rect 577256 421024 578882 421260
rect 490482 420788 578882 421024
rect 490482 420552 572772 420788
rect 573008 420552 573244 420788
rect 573480 420552 573716 420788
rect 573952 420552 574188 420788
rect 574424 420552 574660 420788
rect 574896 420552 575132 420788
rect 575368 420552 575604 420788
rect 575840 420552 576076 420788
rect 576312 420552 576548 420788
rect 576784 420552 577020 420788
rect 577256 420552 578882 420788
rect -800 420358 480 420470
rect 490482 420272 578882 420552
rect -800 419176 480 419288
rect 583520 411206 584800 411318
rect 583520 410024 584800 410136
rect 583520 408842 584800 408954
rect 583520 407660 584800 407772
rect 583520 406478 584800 406590
rect 583520 405296 584800 405408
rect -800 381864 480 381976
rect -800 380682 480 380794
rect -800 379500 480 379612
rect -800 378318 480 378430
rect 477192 377866 483800 378072
rect 477060 377836 567660 377866
rect 477060 377600 477192 377836
rect 477428 377600 477664 377836
rect 477900 377600 478136 377836
rect 478372 377600 478608 377836
rect 478844 377600 479080 377836
rect 479316 377600 479552 377836
rect 479788 377600 480024 377836
rect 480260 377600 480496 377836
rect 480732 377600 480968 377836
rect 481204 377600 481440 377836
rect 481676 377600 481912 377836
rect 482148 377600 482384 377836
rect 482620 377600 482856 377836
rect 483092 377600 483328 377836
rect 483564 377600 567660 377836
rect 477060 377364 562624 377600
rect 562860 377364 563096 377600
rect 563332 377364 563568 377600
rect 563804 377364 564040 377600
rect 564276 377364 564512 377600
rect 564748 377364 564984 377600
rect 565220 377364 565456 377600
rect 565692 377364 565928 377600
rect 566164 377364 566400 377600
rect 566636 377364 566872 377600
rect 567108 377364 567660 377600
rect -800 377136 480 377248
rect 477060 377128 477192 377364
rect 477428 377128 477664 377364
rect 477900 377128 478136 377364
rect 478372 377128 478608 377364
rect 478844 377128 479080 377364
rect 479316 377128 479552 377364
rect 479788 377128 480024 377364
rect 480260 377128 480496 377364
rect 480732 377128 480968 377364
rect 481204 377128 481440 377364
rect 481676 377128 481912 377364
rect 482148 377128 482384 377364
rect 482620 377128 482856 377364
rect 483092 377128 483328 377364
rect 483564 377128 567660 377364
rect 477060 376892 562624 377128
rect 562860 376892 563096 377128
rect 563332 376892 563568 377128
rect 563804 376892 564040 377128
rect 564276 376892 564512 377128
rect 564748 376892 564984 377128
rect 565220 376892 565456 377128
rect 565692 376892 565928 377128
rect 566164 376892 566400 377128
rect 566636 376892 566872 377128
rect 567108 376892 567660 377128
rect 477060 376656 477192 376892
rect 477428 376656 477664 376892
rect 477900 376656 478136 376892
rect 478372 376656 478608 376892
rect 478844 376656 479080 376892
rect 479316 376656 479552 376892
rect 479788 376656 480024 376892
rect 480260 376656 480496 376892
rect 480732 376656 480968 376892
rect 481204 376656 481440 376892
rect 481676 376656 481912 376892
rect 482148 376656 482384 376892
rect 482620 376656 482856 376892
rect 483092 376656 483328 376892
rect 483564 376656 567660 376892
rect 477060 376420 562624 376656
rect 562860 376420 563096 376656
rect 563332 376420 563568 376656
rect 563804 376420 564040 376656
rect 564276 376420 564512 376656
rect 564748 376420 564984 376656
rect 565220 376420 565456 376656
rect 565692 376420 565928 376656
rect 566164 376420 566400 376656
rect 566636 376420 566872 376656
rect 567108 376420 567660 376656
rect 477060 376184 477192 376420
rect 477428 376184 477664 376420
rect 477900 376184 478136 376420
rect 478372 376184 478608 376420
rect 478844 376184 479080 376420
rect 479316 376184 479552 376420
rect 479788 376184 480024 376420
rect 480260 376184 480496 376420
rect 480732 376184 480968 376420
rect 481204 376184 481440 376420
rect 481676 376184 481912 376420
rect 482148 376184 482384 376420
rect 482620 376184 482856 376420
rect 483092 376184 483328 376420
rect 483564 376184 567660 376420
rect -800 375954 480 376066
rect 477060 375948 562624 376184
rect 562860 375948 563096 376184
rect 563332 375948 563568 376184
rect 563804 375948 564040 376184
rect 564276 375948 564512 376184
rect 564748 375948 564984 376184
rect 565220 375948 565456 376184
rect 565692 375948 565928 376184
rect 566164 375948 566400 376184
rect 566636 375948 566872 376184
rect 567108 375948 567660 376184
rect 477060 375712 477192 375948
rect 477428 375712 477664 375948
rect 477900 375712 478136 375948
rect 478372 375712 478608 375948
rect 478844 375712 479080 375948
rect 479316 375712 479552 375948
rect 479788 375712 480024 375948
rect 480260 375712 480496 375948
rect 480732 375712 480968 375948
rect 481204 375712 481440 375948
rect 481676 375712 481912 375948
rect 482148 375712 482384 375948
rect 482620 375712 482856 375948
rect 483092 375712 483328 375948
rect 483564 375712 567660 375948
rect 477060 375476 562624 375712
rect 562860 375476 563096 375712
rect 563332 375476 563568 375712
rect 563804 375476 564040 375712
rect 564276 375476 564512 375712
rect 564748 375476 564984 375712
rect 565220 375476 565456 375712
rect 565692 375476 565928 375712
rect 566164 375476 566400 375712
rect 566636 375476 566872 375712
rect 567108 375476 567660 375712
rect 477060 375240 477192 375476
rect 477428 375240 477664 375476
rect 477900 375240 478136 375476
rect 478372 375240 478608 375476
rect 478844 375240 479080 375476
rect 479316 375240 479552 375476
rect 479788 375240 480024 375476
rect 480260 375240 480496 375476
rect 480732 375240 480968 375476
rect 481204 375240 481440 375476
rect 481676 375240 481912 375476
rect 482148 375240 482384 375476
rect 482620 375240 482856 375476
rect 483092 375240 483328 375476
rect 483564 375240 567660 375476
rect 477060 375004 562624 375240
rect 562860 375004 563096 375240
rect 563332 375004 563568 375240
rect 563804 375004 564040 375240
rect 564276 375004 564512 375240
rect 564748 375004 564984 375240
rect 565220 375004 565456 375240
rect 565692 375004 565928 375240
rect 566164 375004 566400 375240
rect 566636 375004 566872 375240
rect 567108 375004 567660 375240
rect 477060 374768 477192 375004
rect 477428 374768 477664 375004
rect 477900 374768 478136 375004
rect 478372 374768 478608 375004
rect 478844 374768 479080 375004
rect 479316 374768 479552 375004
rect 479788 374768 480024 375004
rect 480260 374768 480496 375004
rect 480732 374768 480968 375004
rect 481204 374768 481440 375004
rect 481676 374768 481912 375004
rect 482148 374768 482384 375004
rect 482620 374768 482856 375004
rect 483092 374768 483328 375004
rect 483564 374768 567660 375004
rect 477060 374532 562624 374768
rect 562860 374532 563096 374768
rect 563332 374532 563568 374768
rect 563804 374532 564040 374768
rect 564276 374532 564512 374768
rect 564748 374532 564984 374768
rect 565220 374532 565456 374768
rect 565692 374532 565928 374768
rect 566164 374532 566400 374768
rect 566636 374532 566872 374768
rect 567108 374532 567660 374768
rect 477060 374296 477192 374532
rect 477428 374296 477664 374532
rect 477900 374296 478136 374532
rect 478372 374296 478608 374532
rect 478844 374296 479080 374532
rect 479316 374296 479552 374532
rect 479788 374296 480024 374532
rect 480260 374296 480496 374532
rect 480732 374296 480968 374532
rect 481204 374296 481440 374532
rect 481676 374296 481912 374532
rect 482148 374296 482384 374532
rect 482620 374296 482856 374532
rect 483092 374296 483328 374532
rect 483564 374296 567660 374532
rect 477060 374060 562624 374296
rect 562860 374060 563096 374296
rect 563332 374060 563568 374296
rect 563804 374060 564040 374296
rect 564276 374060 564512 374296
rect 564748 374060 564984 374296
rect 565220 374060 565456 374296
rect 565692 374060 565928 374296
rect 566164 374060 566400 374296
rect 566636 374060 566872 374296
rect 567108 374060 567660 374296
rect 477060 373824 477192 374060
rect 477428 373824 477664 374060
rect 477900 373824 478136 374060
rect 478372 373824 478608 374060
rect 478844 373824 479080 374060
rect 479316 373824 479552 374060
rect 479788 373824 480024 374060
rect 480260 373824 480496 374060
rect 480732 373824 480968 374060
rect 481204 373824 481440 374060
rect 481676 373824 481912 374060
rect 482148 373824 482384 374060
rect 482620 373824 482856 374060
rect 483092 373824 483328 374060
rect 483564 373824 567660 374060
rect 477060 373588 562624 373824
rect 562860 373588 563096 373824
rect 563332 373588 563568 373824
rect 563804 373588 564040 373824
rect 564276 373588 564512 373824
rect 564748 373588 564984 373824
rect 565220 373588 565456 373824
rect 565692 373588 565928 373824
rect 566164 373588 566400 373824
rect 566636 373588 566872 373824
rect 567108 373588 567660 373824
rect 477060 373352 477192 373588
rect 477428 373352 477664 373588
rect 477900 373352 478136 373588
rect 478372 373352 478608 373588
rect 478844 373352 479080 373588
rect 479316 373352 479552 373588
rect 479788 373352 480024 373588
rect 480260 373352 480496 373588
rect 480732 373352 480968 373588
rect 481204 373352 481440 373588
rect 481676 373352 481912 373588
rect 482148 373352 482384 373588
rect 482620 373352 482856 373588
rect 483092 373352 483328 373588
rect 483564 373352 567660 373588
rect 477060 373116 562624 373352
rect 562860 373116 563096 373352
rect 563332 373116 563568 373352
rect 563804 373116 564040 373352
rect 564276 373116 564512 373352
rect 564748 373116 564984 373352
rect 565220 373116 565456 373352
rect 565692 373116 565928 373352
rect 566164 373116 566400 373352
rect 566636 373116 566872 373352
rect 567108 373116 567660 373352
rect 477060 372880 477192 373116
rect 477428 372880 477664 373116
rect 477900 372880 478136 373116
rect 478372 372880 478608 373116
rect 478844 372880 479080 373116
rect 479316 372880 479552 373116
rect 479788 372880 480024 373116
rect 480260 372880 480496 373116
rect 480732 372880 480968 373116
rect 481204 372880 481440 373116
rect 481676 372880 481912 373116
rect 482148 372880 482384 373116
rect 482620 372880 482856 373116
rect 483092 372880 483328 373116
rect 483564 372880 567660 373116
rect 477060 372644 562624 372880
rect 562860 372644 563096 372880
rect 563332 372644 563568 372880
rect 563804 372644 564040 372880
rect 564276 372644 564512 372880
rect 564748 372644 564984 372880
rect 565220 372644 565456 372880
rect 565692 372644 565928 372880
rect 566164 372644 566400 372880
rect 566636 372644 566872 372880
rect 567108 372644 567660 372880
rect 477060 372408 477192 372644
rect 477428 372408 477664 372644
rect 477900 372408 478136 372644
rect 478372 372408 478608 372644
rect 478844 372408 479080 372644
rect 479316 372408 479552 372644
rect 479788 372408 480024 372644
rect 480260 372408 480496 372644
rect 480732 372408 480968 372644
rect 481204 372408 481440 372644
rect 481676 372408 481912 372644
rect 482148 372408 482384 372644
rect 482620 372408 482856 372644
rect 483092 372408 483328 372644
rect 483564 372408 567660 372644
rect 477060 372172 562624 372408
rect 562860 372172 563096 372408
rect 563332 372172 563568 372408
rect 563804 372172 564040 372408
rect 564276 372172 564512 372408
rect 564748 372172 564984 372408
rect 565220 372172 565456 372408
rect 565692 372172 565928 372408
rect 566164 372172 566400 372408
rect 566636 372172 566872 372408
rect 567108 372172 567660 372408
rect 477060 371936 477192 372172
rect 477428 371936 477664 372172
rect 477900 371936 478136 372172
rect 478372 371936 478608 372172
rect 478844 371936 479080 372172
rect 479316 371936 479552 372172
rect 479788 371936 480024 372172
rect 480260 371936 480496 372172
rect 480732 371936 480968 372172
rect 481204 371936 481440 372172
rect 481676 371936 481912 372172
rect 482148 371936 482384 372172
rect 482620 371936 482856 372172
rect 483092 371936 483328 372172
rect 483564 371936 567660 372172
rect 477060 371700 562624 371936
rect 562860 371700 563096 371936
rect 563332 371700 563568 371936
rect 563804 371700 564040 371936
rect 564276 371700 564512 371936
rect 564748 371700 564984 371936
rect 565220 371700 565456 371936
rect 565692 371700 565928 371936
rect 566164 371700 566400 371936
rect 566636 371700 566872 371936
rect 567108 371700 567660 371936
rect 477060 371464 477192 371700
rect 477428 371464 477664 371700
rect 477900 371464 478136 371700
rect 478372 371464 478608 371700
rect 478844 371464 479080 371700
rect 479316 371464 479552 371700
rect 479788 371464 480024 371700
rect 480260 371464 480496 371700
rect 480732 371464 480968 371700
rect 481204 371464 481440 371700
rect 481676 371464 481912 371700
rect 482148 371464 482384 371700
rect 482620 371464 482856 371700
rect 483092 371464 483328 371700
rect 483564 371464 567660 371700
rect 477060 371228 562624 371464
rect 562860 371228 563096 371464
rect 563332 371228 563568 371464
rect 563804 371228 564040 371464
rect 564276 371228 564512 371464
rect 564748 371228 564984 371464
rect 565220 371228 565456 371464
rect 565692 371228 565928 371464
rect 566164 371228 566400 371464
rect 566636 371228 566872 371464
rect 567108 371228 567660 371464
rect 477060 371200 567660 371228
rect 583520 364784 584800 364896
rect 583520 363602 584800 363714
rect 583520 362420 584800 362532
rect 583520 361238 584800 361350
rect 583520 360056 584800 360168
rect 583520 358874 584800 358986
rect -800 338642 480 338754
rect -800 337460 480 337572
rect -800 336278 480 336390
rect -800 335096 480 335208
rect -800 333914 480 334026
rect -800 332732 480 332844
rect 583520 319562 584800 319674
rect 583520 318380 584800 318492
rect 583520 317198 584800 317310
rect 583520 316016 584800 316128
rect 583520 314834 584800 314946
rect 583520 313652 584800 313764
rect -800 295420 480 295532
rect -800 294238 480 294350
rect -800 293056 480 293168
rect -800 291874 480 291986
rect -800 290692 480 290804
rect -800 289510 480 289622
rect 583520 275140 584800 275252
rect 583520 273958 584800 274070
rect 583520 272776 584800 272888
rect 583520 271594 584800 271706
rect 583520 270412 584800 270524
rect 583520 269230 584800 269342
rect -800 252398 480 252510
rect -800 251216 480 251328
rect -800 250034 480 250146
rect -800 248852 480 248964
rect -800 247670 480 247782
rect -800 246488 480 246600
rect 582340 235230 584800 240030
rect 582340 225230 584800 230030
rect -800 214888 1660 219688
rect -800 204888 1660 209688
rect 582340 191430 584800 196230
rect 582340 181430 584800 186230
rect -800 172888 1660 177688
rect -800 162888 1660 167688
rect 582340 146830 584800 151630
rect 582340 136830 584800 141630
rect -800 124776 480 124888
rect -800 123594 480 123706
rect -800 122412 480 122524
rect -800 121230 480 121342
rect -800 120048 480 120160
rect -800 118866 480 118978
rect 583520 95118 584800 95230
rect 583520 93936 584800 94048
rect 583520 92754 584800 92866
rect 583520 91572 584800 91684
rect -800 81554 480 81666
rect -800 80372 480 80484
rect -800 79190 480 79302
rect -800 78008 480 78120
rect -800 76826 480 76938
rect -800 75644 480 75756
rect 583520 50460 584800 50572
rect 583520 49278 584800 49390
rect 583520 48096 584800 48208
rect 583520 46914 584800 47026
rect -800 38332 480 38444
rect -800 37150 480 37262
rect -800 35968 480 36080
rect -800 34786 480 34898
rect -800 33604 480 33716
rect -800 32422 480 32534
rect 583520 24002 584800 24114
rect 583520 22820 584800 22932
rect 583520 21638 584800 21750
rect 583520 20456 584800 20568
rect 583520 19274 584800 19386
rect 583520 18092 584800 18204
rect -800 16910 480 17022
rect 583520 16910 584800 17022
rect -800 15728 480 15840
rect 583520 15728 584800 15840
rect -800 14546 480 14658
rect 583520 14546 584800 14658
rect -800 13364 480 13476
rect 583520 13364 584800 13476
rect -800 12182 480 12294
rect 583520 12182 584800 12294
rect -800 11000 480 11112
rect 583520 11000 584800 11112
rect -800 9818 480 9930
rect 583520 9818 584800 9930
rect -800 8636 480 8748
rect 583520 8636 584800 8748
rect -800 7454 480 7566
rect 583520 7454 584800 7566
rect -800 6272 480 6384
rect 583520 6272 584800 6384
rect -800 5090 480 5202
rect 583520 5090 584800 5202
rect -800 3908 480 4020
rect 583520 3908 584800 4020
rect -800 2726 480 2838
rect 583520 2726 584800 2838
rect -800 1544 480 1656
rect 583520 1544 584800 1656
<< via3 >>
rect 171000 692600 173000 697200
rect 173400 692600 175400 697200
rect 222706 692600 224706 697200
rect 225106 692600 227106 697200
rect 324412 692600 326412 697200
rect 326812 692600 328812 697200
rect 510654 692560 515334 697360
rect 520654 692560 525334 697360
rect 562600 639844 567400 644524
rect 562600 629844 567400 634524
rect 477192 522626 477428 522862
rect 477664 522626 477900 522862
rect 478136 522626 478372 522862
rect 478608 522626 478844 522862
rect 479080 522626 479316 522862
rect 479552 522626 479788 522862
rect 480024 522626 480260 522862
rect 480496 522626 480732 522862
rect 480968 522626 481204 522862
rect 481440 522626 481676 522862
rect 481912 522626 482148 522862
rect 482384 522626 482620 522862
rect 482856 522626 483092 522862
rect 483328 522626 483564 522862
rect 562624 522504 562860 522740
rect 563096 522504 563332 522740
rect 563568 522504 563804 522740
rect 564040 522504 564276 522740
rect 564512 522504 564748 522740
rect 564984 522504 565220 522740
rect 565456 522504 565692 522740
rect 565928 522504 566164 522740
rect 566400 522504 566636 522740
rect 566872 522504 567108 522740
rect 477192 522154 477428 522390
rect 477664 522154 477900 522390
rect 478136 522154 478372 522390
rect 478608 522154 478844 522390
rect 479080 522154 479316 522390
rect 479552 522154 479788 522390
rect 480024 522154 480260 522390
rect 480496 522154 480732 522390
rect 480968 522154 481204 522390
rect 481440 522154 481676 522390
rect 481912 522154 482148 522390
rect 482384 522154 482620 522390
rect 482856 522154 483092 522390
rect 483328 522154 483564 522390
rect 562624 522032 562860 522268
rect 563096 522032 563332 522268
rect 563568 522032 563804 522268
rect 564040 522032 564276 522268
rect 564512 522032 564748 522268
rect 564984 522032 565220 522268
rect 565456 522032 565692 522268
rect 565928 522032 566164 522268
rect 566400 522032 566636 522268
rect 566872 522032 567108 522268
rect 477192 521682 477428 521918
rect 477664 521682 477900 521918
rect 478136 521682 478372 521918
rect 478608 521682 478844 521918
rect 479080 521682 479316 521918
rect 479552 521682 479788 521918
rect 480024 521682 480260 521918
rect 480496 521682 480732 521918
rect 480968 521682 481204 521918
rect 481440 521682 481676 521918
rect 481912 521682 482148 521918
rect 482384 521682 482620 521918
rect 482856 521682 483092 521918
rect 483328 521682 483564 521918
rect 562624 521560 562860 521796
rect 563096 521560 563332 521796
rect 563568 521560 563804 521796
rect 564040 521560 564276 521796
rect 564512 521560 564748 521796
rect 564984 521560 565220 521796
rect 565456 521560 565692 521796
rect 565928 521560 566164 521796
rect 566400 521560 566636 521796
rect 566872 521560 567108 521796
rect 477192 521210 477428 521446
rect 477664 521210 477900 521446
rect 478136 521210 478372 521446
rect 478608 521210 478844 521446
rect 479080 521210 479316 521446
rect 479552 521210 479788 521446
rect 480024 521210 480260 521446
rect 480496 521210 480732 521446
rect 480968 521210 481204 521446
rect 481440 521210 481676 521446
rect 481912 521210 482148 521446
rect 482384 521210 482620 521446
rect 482856 521210 483092 521446
rect 483328 521210 483564 521446
rect 562624 521088 562860 521324
rect 563096 521088 563332 521324
rect 563568 521088 563804 521324
rect 564040 521088 564276 521324
rect 564512 521088 564748 521324
rect 564984 521088 565220 521324
rect 565456 521088 565692 521324
rect 565928 521088 566164 521324
rect 566400 521088 566636 521324
rect 566872 521088 567108 521324
rect 477192 520738 477428 520974
rect 477664 520738 477900 520974
rect 478136 520738 478372 520974
rect 478608 520738 478844 520974
rect 479080 520738 479316 520974
rect 479552 520738 479788 520974
rect 480024 520738 480260 520974
rect 480496 520738 480732 520974
rect 480968 520738 481204 520974
rect 481440 520738 481676 520974
rect 481912 520738 482148 520974
rect 482384 520738 482620 520974
rect 482856 520738 483092 520974
rect 483328 520738 483564 520974
rect 562624 520616 562860 520852
rect 563096 520616 563332 520852
rect 563568 520616 563804 520852
rect 564040 520616 564276 520852
rect 564512 520616 564748 520852
rect 564984 520616 565220 520852
rect 565456 520616 565692 520852
rect 565928 520616 566164 520852
rect 566400 520616 566636 520852
rect 566872 520616 567108 520852
rect 477192 520266 477428 520502
rect 477664 520266 477900 520502
rect 478136 520266 478372 520502
rect 478608 520266 478844 520502
rect 479080 520266 479316 520502
rect 479552 520266 479788 520502
rect 480024 520266 480260 520502
rect 480496 520266 480732 520502
rect 480968 520266 481204 520502
rect 481440 520266 481676 520502
rect 481912 520266 482148 520502
rect 482384 520266 482620 520502
rect 482856 520266 483092 520502
rect 483328 520266 483564 520502
rect 562624 520144 562860 520380
rect 563096 520144 563332 520380
rect 563568 520144 563804 520380
rect 564040 520144 564276 520380
rect 564512 520144 564748 520380
rect 564984 520144 565220 520380
rect 565456 520144 565692 520380
rect 565928 520144 566164 520380
rect 566400 520144 566636 520380
rect 566872 520144 567108 520380
rect 477192 519794 477428 520030
rect 477664 519794 477900 520030
rect 478136 519794 478372 520030
rect 478608 519794 478844 520030
rect 479080 519794 479316 520030
rect 479552 519794 479788 520030
rect 480024 519794 480260 520030
rect 480496 519794 480732 520030
rect 480968 519794 481204 520030
rect 481440 519794 481676 520030
rect 481912 519794 482148 520030
rect 482384 519794 482620 520030
rect 482856 519794 483092 520030
rect 483328 519794 483564 520030
rect 562624 519672 562860 519908
rect 563096 519672 563332 519908
rect 563568 519672 563804 519908
rect 564040 519672 564276 519908
rect 564512 519672 564748 519908
rect 564984 519672 565220 519908
rect 565456 519672 565692 519908
rect 565928 519672 566164 519908
rect 566400 519672 566636 519908
rect 566872 519672 567108 519908
rect 477192 519322 477428 519558
rect 477664 519322 477900 519558
rect 478136 519322 478372 519558
rect 478608 519322 478844 519558
rect 479080 519322 479316 519558
rect 479552 519322 479788 519558
rect 480024 519322 480260 519558
rect 480496 519322 480732 519558
rect 480968 519322 481204 519558
rect 481440 519322 481676 519558
rect 481912 519322 482148 519558
rect 482384 519322 482620 519558
rect 482856 519322 483092 519558
rect 483328 519322 483564 519558
rect 562624 519200 562860 519436
rect 563096 519200 563332 519436
rect 563568 519200 563804 519436
rect 564040 519200 564276 519436
rect 564512 519200 564748 519436
rect 564984 519200 565220 519436
rect 565456 519200 565692 519436
rect 565928 519200 566164 519436
rect 566400 519200 566636 519436
rect 566872 519200 567108 519436
rect 477192 518850 477428 519086
rect 477664 518850 477900 519086
rect 478136 518850 478372 519086
rect 478608 518850 478844 519086
rect 479080 518850 479316 519086
rect 479552 518850 479788 519086
rect 480024 518850 480260 519086
rect 480496 518850 480732 519086
rect 480968 518850 481204 519086
rect 481440 518850 481676 519086
rect 481912 518850 482148 519086
rect 482384 518850 482620 519086
rect 482856 518850 483092 519086
rect 483328 518850 483564 519086
rect 562624 518728 562860 518964
rect 563096 518728 563332 518964
rect 563568 518728 563804 518964
rect 564040 518728 564276 518964
rect 564512 518728 564748 518964
rect 564984 518728 565220 518964
rect 565456 518728 565692 518964
rect 565928 518728 566164 518964
rect 566400 518728 566636 518964
rect 566872 518728 567108 518964
rect 477192 518378 477428 518614
rect 477664 518378 477900 518614
rect 478136 518378 478372 518614
rect 478608 518378 478844 518614
rect 479080 518378 479316 518614
rect 479552 518378 479788 518614
rect 480024 518378 480260 518614
rect 480496 518378 480732 518614
rect 480968 518378 481204 518614
rect 481440 518378 481676 518614
rect 481912 518378 482148 518614
rect 482384 518378 482620 518614
rect 482856 518378 483092 518614
rect 483328 518378 483564 518614
rect 562624 518256 562860 518492
rect 563096 518256 563332 518492
rect 563568 518256 563804 518492
rect 564040 518256 564276 518492
rect 564512 518256 564748 518492
rect 564984 518256 565220 518492
rect 565456 518256 565692 518492
rect 565928 518256 566164 518492
rect 566400 518256 566636 518492
rect 566872 518256 567108 518492
rect 477192 517906 477428 518142
rect 477664 517906 477900 518142
rect 478136 517906 478372 518142
rect 478608 517906 478844 518142
rect 479080 517906 479316 518142
rect 479552 517906 479788 518142
rect 480024 517906 480260 518142
rect 480496 517906 480732 518142
rect 480968 517906 481204 518142
rect 481440 517906 481676 518142
rect 481912 517906 482148 518142
rect 482384 517906 482620 518142
rect 482856 517906 483092 518142
rect 483328 517906 483564 518142
rect 562624 517784 562860 518020
rect 563096 517784 563332 518020
rect 563568 517784 563804 518020
rect 564040 517784 564276 518020
rect 564512 517784 564748 518020
rect 564984 517784 565220 518020
rect 565456 517784 565692 518020
rect 565928 517784 566164 518020
rect 566400 517784 566636 518020
rect 566872 517784 567108 518020
rect 477192 517434 477428 517670
rect 477664 517434 477900 517670
rect 478136 517434 478372 517670
rect 478608 517434 478844 517670
rect 479080 517434 479316 517670
rect 479552 517434 479788 517670
rect 480024 517434 480260 517670
rect 480496 517434 480732 517670
rect 480968 517434 481204 517670
rect 481440 517434 481676 517670
rect 481912 517434 482148 517670
rect 482384 517434 482620 517670
rect 482856 517434 483092 517670
rect 483328 517434 483564 517670
rect 562624 517312 562860 517548
rect 563096 517312 563332 517548
rect 563568 517312 563804 517548
rect 564040 517312 564276 517548
rect 564512 517312 564748 517548
rect 564984 517312 565220 517548
rect 565456 517312 565692 517548
rect 565928 517312 566164 517548
rect 566400 517312 566636 517548
rect 566872 517312 567108 517548
rect 477192 516962 477428 517198
rect 477664 516962 477900 517198
rect 478136 516962 478372 517198
rect 478608 516962 478844 517198
rect 479080 516962 479316 517198
rect 479552 516962 479788 517198
rect 480024 516962 480260 517198
rect 480496 516962 480732 517198
rect 480968 516962 481204 517198
rect 481440 516962 481676 517198
rect 481912 516962 482148 517198
rect 482384 516962 482620 517198
rect 482856 516962 483092 517198
rect 483328 516962 483564 517198
rect 562624 516840 562860 517076
rect 563096 516840 563332 517076
rect 563568 516840 563804 517076
rect 564040 516840 564276 517076
rect 564512 516840 564748 517076
rect 564984 516840 565220 517076
rect 565456 516840 565692 517076
rect 565928 516840 566164 517076
rect 566400 516840 566636 517076
rect 566872 516840 567108 517076
rect 477192 516490 477428 516726
rect 477664 516490 477900 516726
rect 478136 516490 478372 516726
rect 478608 516490 478844 516726
rect 479080 516490 479316 516726
rect 479552 516490 479788 516726
rect 480024 516490 480260 516726
rect 480496 516490 480732 516726
rect 480968 516490 481204 516726
rect 481440 516490 481676 516726
rect 481912 516490 482148 516726
rect 482384 516490 482620 516726
rect 482856 516490 483092 516726
rect 483328 516490 483564 516726
rect 562624 516368 562860 516604
rect 563096 516368 563332 516604
rect 563568 516368 563804 516604
rect 564040 516368 564276 516604
rect 564512 516368 564748 516604
rect 564984 516368 565220 516604
rect 565456 516368 565692 516604
rect 565928 516368 566164 516604
rect 566400 516368 566636 516604
rect 566872 516368 567108 516604
rect 562480 495662 562560 495742
rect 562640 495662 562720 495742
rect 562800 495662 562880 495742
rect 562960 495662 563040 495742
rect 563120 495662 563200 495742
rect 563280 495662 563360 495742
rect 563440 495662 563520 495742
rect 563600 495662 563680 495742
rect 563760 495662 563840 495742
rect 563920 495662 564000 495742
rect 564080 495662 564160 495742
rect 564240 495662 564320 495742
rect 564400 495662 564480 495742
rect 564560 495662 564640 495742
rect 564720 495662 564800 495742
rect 564880 495662 564960 495742
rect 565040 495662 565120 495742
rect 565200 495662 565280 495742
rect 565360 495662 565440 495742
rect 565520 495662 565600 495742
rect 565680 495662 565760 495742
rect 565840 495662 565920 495742
rect 566000 495662 566080 495742
rect 566160 495662 566240 495742
rect 566320 495662 566400 495742
rect 566480 495662 566560 495742
rect 566640 495662 566720 495742
rect 566800 495662 566880 495742
rect 566960 495662 567040 495742
rect 567120 495662 567200 495742
rect 567280 495662 567360 495742
rect 562480 495502 562560 495582
rect 562640 495502 562720 495582
rect 562800 495502 562880 495582
rect 562960 495502 563040 495582
rect 563120 495502 563200 495582
rect 563280 495502 563360 495582
rect 563440 495502 563520 495582
rect 563600 495502 563680 495582
rect 563760 495502 563840 495582
rect 563920 495502 564000 495582
rect 564080 495502 564160 495582
rect 564240 495502 564320 495582
rect 564400 495502 564480 495582
rect 564560 495502 564640 495582
rect 564720 495502 564800 495582
rect 564880 495502 564960 495582
rect 565040 495502 565120 495582
rect 565200 495502 565280 495582
rect 565360 495502 565440 495582
rect 565520 495502 565600 495582
rect 565680 495502 565760 495582
rect 565840 495502 565920 495582
rect 566000 495502 566080 495582
rect 566160 495502 566240 495582
rect 566320 495502 566400 495582
rect 566480 495502 566560 495582
rect 566640 495502 566720 495582
rect 566800 495502 566880 495582
rect 566960 495502 567040 495582
rect 567120 495502 567200 495582
rect 567280 495502 567360 495582
rect 572640 495662 572720 495742
rect 572800 495662 572880 495742
rect 572960 495662 573040 495742
rect 573120 495662 573200 495742
rect 573280 495662 573360 495742
rect 573440 495662 573520 495742
rect 573600 495662 573680 495742
rect 573760 495662 573840 495742
rect 573920 495662 574000 495742
rect 574080 495662 574160 495742
rect 574240 495662 574320 495742
rect 574400 495662 574480 495742
rect 574560 495662 574640 495742
rect 574720 495662 574800 495742
rect 574880 495662 574960 495742
rect 575040 495662 575120 495742
rect 575200 495662 575280 495742
rect 575360 495662 575440 495742
rect 575520 495662 575600 495742
rect 575680 495662 575760 495742
rect 575840 495662 575920 495742
rect 576000 495662 576080 495742
rect 576160 495662 576240 495742
rect 576320 495662 576400 495742
rect 576480 495662 576560 495742
rect 576640 495662 576720 495742
rect 576800 495662 576880 495742
rect 576960 495662 577040 495742
rect 577120 495662 577200 495742
rect 577280 495662 577360 495742
rect 577440 495662 577520 495742
rect 572640 495502 572720 495582
rect 572800 495502 572880 495582
rect 572960 495502 573040 495582
rect 573120 495502 573200 495582
rect 573280 495502 573360 495582
rect 573440 495502 573520 495582
rect 573600 495502 573680 495582
rect 573760 495502 573840 495582
rect 573920 495502 574000 495582
rect 574080 495502 574160 495582
rect 574240 495502 574320 495582
rect 574400 495502 574480 495582
rect 574560 495502 574640 495582
rect 574720 495502 574800 495582
rect 574880 495502 574960 495582
rect 575040 495502 575120 495582
rect 575200 495502 575280 495582
rect 575360 495502 575440 495582
rect 575520 495502 575600 495582
rect 575680 495502 575760 495582
rect 575840 495502 575920 495582
rect 576000 495502 576080 495582
rect 576160 495502 576240 495582
rect 576320 495502 576400 495582
rect 576480 495502 576560 495582
rect 576640 495502 576720 495582
rect 576800 495502 576880 495582
rect 576960 495502 577040 495582
rect 577120 495502 577200 495582
rect 577280 495502 577360 495582
rect 577440 495502 577520 495582
rect 511616 494464 511680 494528
rect 511744 494464 511808 494528
rect 511872 494464 511936 494528
rect 512000 494464 512064 494528
rect 511616 494336 511680 494400
rect 511744 494336 511808 494400
rect 511872 494336 511936 494400
rect 512000 494336 512064 494400
rect 511616 494208 511680 494272
rect 511744 494208 511808 494272
rect 511872 494208 511936 494272
rect 512000 494208 512064 494272
rect 511616 494080 511680 494144
rect 511744 494080 511808 494144
rect 511872 494080 511936 494144
rect 512000 494080 512064 494144
rect 511616 493952 511680 494016
rect 511744 493952 511808 494016
rect 511872 493952 511936 494016
rect 512000 493952 512064 494016
rect 511616 493824 511680 493888
rect 511744 493824 511808 493888
rect 511872 493824 511936 493888
rect 512000 493824 512064 493888
rect 572772 483564 573008 483800
rect 573244 483564 573480 483800
rect 573716 483564 573952 483800
rect 574188 483564 574424 483800
rect 574660 483564 574896 483800
rect 575132 483564 575368 483800
rect 575604 483564 575840 483800
rect 576076 483564 576312 483800
rect 576548 483564 576784 483800
rect 577020 483564 577256 483800
rect 490940 478452 496684 483236
rect 503960 478452 509704 483236
rect 517360 478452 523104 483236
rect 530760 478452 536504 483236
rect 572772 483092 573008 483328
rect 573244 483092 573480 483328
rect 573716 483092 573952 483328
rect 574188 483092 574424 483328
rect 574660 483092 574896 483328
rect 575132 483092 575368 483328
rect 575604 483092 575840 483328
rect 576076 483092 576312 483328
rect 576548 483092 576784 483328
rect 577020 483092 577256 483328
rect 572772 482620 573008 482856
rect 573244 482620 573480 482856
rect 573716 482620 573952 482856
rect 574188 482620 574424 482856
rect 574660 482620 574896 482856
rect 575132 482620 575368 482856
rect 575604 482620 575840 482856
rect 576076 482620 576312 482856
rect 576548 482620 576784 482856
rect 577020 482620 577256 482856
rect 572772 482148 573008 482384
rect 573244 482148 573480 482384
rect 573716 482148 573952 482384
rect 574188 482148 574424 482384
rect 574660 482148 574896 482384
rect 575132 482148 575368 482384
rect 575604 482148 575840 482384
rect 576076 482148 576312 482384
rect 576548 482148 576784 482384
rect 577020 482148 577256 482384
rect 572772 481676 573008 481912
rect 573244 481676 573480 481912
rect 573716 481676 573952 481912
rect 574188 481676 574424 481912
rect 574660 481676 574896 481912
rect 575132 481676 575368 481912
rect 575604 481676 575840 481912
rect 576076 481676 576312 481912
rect 576548 481676 576784 481912
rect 577020 481676 577256 481912
rect 572772 481204 573008 481440
rect 573244 481204 573480 481440
rect 573716 481204 573952 481440
rect 574188 481204 574424 481440
rect 574660 481204 574896 481440
rect 575132 481204 575368 481440
rect 575604 481204 575840 481440
rect 576076 481204 576312 481440
rect 576548 481204 576784 481440
rect 577020 481204 577256 481440
rect 572772 480732 573008 480968
rect 573244 480732 573480 480968
rect 573716 480732 573952 480968
rect 574188 480732 574424 480968
rect 574660 480732 574896 480968
rect 575132 480732 575368 480968
rect 575604 480732 575840 480968
rect 576076 480732 576312 480968
rect 576548 480732 576784 480968
rect 577020 480732 577256 480968
rect 572772 480260 573008 480496
rect 573244 480260 573480 480496
rect 573716 480260 573952 480496
rect 574188 480260 574424 480496
rect 574660 480260 574896 480496
rect 575132 480260 575368 480496
rect 575604 480260 575840 480496
rect 576076 480260 576312 480496
rect 576548 480260 576784 480496
rect 577020 480260 577256 480496
rect 572772 479788 573008 480024
rect 573244 479788 573480 480024
rect 573716 479788 573952 480024
rect 574188 479788 574424 480024
rect 574660 479788 574896 480024
rect 575132 479788 575368 480024
rect 575604 479788 575840 480024
rect 576076 479788 576312 480024
rect 576548 479788 576784 480024
rect 577020 479788 577256 480024
rect 572772 479316 573008 479552
rect 573244 479316 573480 479552
rect 573716 479316 573952 479552
rect 574188 479316 574424 479552
rect 574660 479316 574896 479552
rect 575132 479316 575368 479552
rect 575604 479316 575840 479552
rect 576076 479316 576312 479552
rect 576548 479316 576784 479552
rect 577020 479316 577256 479552
rect 572772 478844 573008 479080
rect 573244 478844 573480 479080
rect 573716 478844 573952 479080
rect 574188 478844 574424 479080
rect 574660 478844 574896 479080
rect 575132 478844 575368 479080
rect 575604 478844 575840 479080
rect 576076 478844 576312 479080
rect 576548 478844 576784 479080
rect 577020 478844 577256 479080
rect 572772 478372 573008 478608
rect 573244 478372 573480 478608
rect 573716 478372 573952 478608
rect 574188 478372 574424 478608
rect 574660 478372 574896 478608
rect 575132 478372 575368 478608
rect 575604 478372 575840 478608
rect 576076 478372 576312 478608
rect 576548 478372 576784 478608
rect 577020 478372 577256 478608
rect 572772 477900 573008 478136
rect 573244 477900 573480 478136
rect 573716 477900 573952 478136
rect 574188 477900 574424 478136
rect 574660 477900 574896 478136
rect 575132 477900 575368 478136
rect 575604 477900 575840 478136
rect 576076 477900 576312 478136
rect 576548 477900 576784 478136
rect 577020 477900 577256 478136
rect 503920 475206 504020 475306
rect 504144 475206 504244 475306
rect 504368 475206 504468 475306
rect 504592 475206 504692 475306
rect 504816 475206 504916 475306
rect 505040 475206 505140 475306
rect 505264 475206 505364 475306
rect 505488 475206 505588 475306
rect 505712 475206 505812 475306
rect 505936 475206 506036 475306
rect 506160 475206 506260 475306
rect 506384 475206 506484 475306
rect 506608 475206 506708 475306
rect 506832 475206 506932 475306
rect 507056 475206 507156 475306
rect 507280 475206 507380 475306
rect 507504 475206 507604 475306
rect 507728 475206 507828 475306
rect 507952 475206 508052 475306
rect 508176 475206 508276 475306
rect 508400 475206 508500 475306
rect 508624 475206 508724 475306
rect 508848 475206 508948 475306
rect 509072 475206 509172 475306
rect 509296 475206 509396 475306
rect 509520 475206 509620 475306
rect 509744 475206 509844 475306
rect 509968 475206 510068 475306
rect 510192 475206 510292 475306
rect 510416 475206 510516 475306
rect 503920 474982 504020 475082
rect 504144 474982 504244 475082
rect 504368 474982 504468 475082
rect 504592 474982 504692 475082
rect 504816 474982 504916 475082
rect 505040 474982 505140 475082
rect 505264 474982 505364 475082
rect 505488 474982 505588 475082
rect 505712 474982 505812 475082
rect 505936 474982 506036 475082
rect 506160 474982 506260 475082
rect 506384 474982 506484 475082
rect 506608 474982 506708 475082
rect 506832 474982 506932 475082
rect 507056 474982 507156 475082
rect 507280 474982 507380 475082
rect 507504 474982 507604 475082
rect 507728 474982 507828 475082
rect 507952 474982 508052 475082
rect 508176 474982 508276 475082
rect 508400 474982 508500 475082
rect 508624 474982 508724 475082
rect 508848 474982 508948 475082
rect 509072 474982 509172 475082
rect 509296 474982 509396 475082
rect 509520 474982 509620 475082
rect 509744 474982 509844 475082
rect 509968 474982 510068 475082
rect 510192 474982 510292 475082
rect 510416 474982 510516 475082
rect 503920 474758 504020 474858
rect 504144 474758 504244 474858
rect 504368 474758 504468 474858
rect 504592 474758 504692 474858
rect 504816 474758 504916 474858
rect 505040 474758 505140 474858
rect 505264 474758 505364 474858
rect 505488 474758 505588 474858
rect 505712 474758 505812 474858
rect 505936 474758 506036 474858
rect 506160 474758 506260 474858
rect 506384 474758 506484 474858
rect 506608 474758 506708 474858
rect 506832 474758 506932 474858
rect 507056 474758 507156 474858
rect 507280 474758 507380 474858
rect 507504 474758 507604 474858
rect 507728 474758 507828 474858
rect 507952 474758 508052 474858
rect 508176 474758 508276 474858
rect 508400 474758 508500 474858
rect 508624 474758 508724 474858
rect 508848 474758 508948 474858
rect 509072 474758 509172 474858
rect 509296 474758 509396 474858
rect 509520 474758 509620 474858
rect 509744 474758 509844 474858
rect 509968 474758 510068 474858
rect 510192 474758 510292 474858
rect 510416 474758 510516 474858
rect 503920 474534 504020 474634
rect 504144 474534 504244 474634
rect 504368 474534 504468 474634
rect 504592 474534 504692 474634
rect 504816 474534 504916 474634
rect 505040 474534 505140 474634
rect 505264 474534 505364 474634
rect 505488 474534 505588 474634
rect 505712 474534 505812 474634
rect 505936 474534 506036 474634
rect 506160 474534 506260 474634
rect 506384 474534 506484 474634
rect 506608 474534 506708 474634
rect 506832 474534 506932 474634
rect 507056 474534 507156 474634
rect 507280 474534 507380 474634
rect 507504 474534 507604 474634
rect 507728 474534 507828 474634
rect 507952 474534 508052 474634
rect 508176 474534 508276 474634
rect 508400 474534 508500 474634
rect 508624 474534 508724 474634
rect 508848 474534 508948 474634
rect 509072 474534 509172 474634
rect 509296 474534 509396 474634
rect 509520 474534 509620 474634
rect 509744 474534 509844 474634
rect 509968 474534 510068 474634
rect 510192 474534 510292 474634
rect 510416 474534 510516 474634
rect 491256 469452 497000 474236
rect 500398 474180 500498 474280
rect 500622 474180 500722 474280
rect 500846 474180 500946 474280
rect 501070 474180 501170 474280
rect 501294 474180 501394 474280
rect 503920 474310 504020 474410
rect 504144 474310 504244 474410
rect 504368 474310 504468 474410
rect 504592 474310 504692 474410
rect 504816 474310 504916 474410
rect 505040 474310 505140 474410
rect 505264 474310 505364 474410
rect 505488 474310 505588 474410
rect 505712 474310 505812 474410
rect 505936 474310 506036 474410
rect 506160 474310 506260 474410
rect 506384 474310 506484 474410
rect 506608 474310 506708 474410
rect 506832 474310 506932 474410
rect 507056 474310 507156 474410
rect 507280 474310 507380 474410
rect 507504 474310 507604 474410
rect 507728 474310 507828 474410
rect 507952 474310 508052 474410
rect 508176 474310 508276 474410
rect 508400 474310 508500 474410
rect 508624 474310 508724 474410
rect 508848 474310 508948 474410
rect 509072 474310 509172 474410
rect 509296 474310 509396 474410
rect 509520 474310 509620 474410
rect 509744 474310 509844 474410
rect 509968 474310 510068 474410
rect 510192 474310 510292 474410
rect 510416 474310 510516 474410
rect 511648 475236 511712 475300
rect 511776 475236 511840 475300
rect 511904 475236 511968 475300
rect 512032 475236 512096 475300
rect 511648 475108 511712 475172
rect 511776 475108 511840 475172
rect 511904 475108 511968 475172
rect 512032 475108 512096 475172
rect 511648 474980 511712 475044
rect 511776 474980 511840 475044
rect 511904 474980 511968 475044
rect 512032 474980 512096 475044
rect 511648 474852 511712 474916
rect 511776 474852 511840 474916
rect 511904 474852 511968 474916
rect 512032 474852 512096 474916
rect 511648 474724 511712 474788
rect 511776 474724 511840 474788
rect 511904 474724 511968 474788
rect 512032 474724 512096 474788
rect 511648 474596 511712 474660
rect 511776 474596 511840 474660
rect 511904 474596 511968 474660
rect 512032 474596 512096 474660
rect 511648 474468 511712 474532
rect 511776 474468 511840 474532
rect 511904 474468 511968 474532
rect 512032 474468 512096 474532
rect 511648 474340 511712 474404
rect 511776 474340 511840 474404
rect 511904 474340 511968 474404
rect 512032 474340 512096 474404
rect 517320 475206 517420 475306
rect 517544 475206 517644 475306
rect 517768 475206 517868 475306
rect 517992 475206 518092 475306
rect 518216 475206 518316 475306
rect 518440 475206 518540 475306
rect 518664 475206 518764 475306
rect 518888 475206 518988 475306
rect 519112 475206 519212 475306
rect 519336 475206 519436 475306
rect 519560 475206 519660 475306
rect 519784 475206 519884 475306
rect 520008 475206 520108 475306
rect 520232 475206 520332 475306
rect 520456 475206 520556 475306
rect 520680 475206 520780 475306
rect 520904 475206 521004 475306
rect 521128 475206 521228 475306
rect 521352 475206 521452 475306
rect 521576 475206 521676 475306
rect 521800 475206 521900 475306
rect 522024 475206 522124 475306
rect 522248 475206 522348 475306
rect 522472 475206 522572 475306
rect 522696 475206 522796 475306
rect 522920 475206 523020 475306
rect 523144 475206 523244 475306
rect 523368 475206 523468 475306
rect 523592 475206 523692 475306
rect 523816 475206 523916 475306
rect 517320 474982 517420 475082
rect 517544 474982 517644 475082
rect 517768 474982 517868 475082
rect 517992 474982 518092 475082
rect 518216 474982 518316 475082
rect 518440 474982 518540 475082
rect 518664 474982 518764 475082
rect 518888 474982 518988 475082
rect 519112 474982 519212 475082
rect 519336 474982 519436 475082
rect 519560 474982 519660 475082
rect 519784 474982 519884 475082
rect 520008 474982 520108 475082
rect 520232 474982 520332 475082
rect 520456 474982 520556 475082
rect 520680 474982 520780 475082
rect 520904 474982 521004 475082
rect 521128 474982 521228 475082
rect 521352 474982 521452 475082
rect 521576 474982 521676 475082
rect 521800 474982 521900 475082
rect 522024 474982 522124 475082
rect 522248 474982 522348 475082
rect 522472 474982 522572 475082
rect 522696 474982 522796 475082
rect 522920 474982 523020 475082
rect 523144 474982 523244 475082
rect 523368 474982 523468 475082
rect 523592 474982 523692 475082
rect 523816 474982 523916 475082
rect 517320 474758 517420 474858
rect 517544 474758 517644 474858
rect 517768 474758 517868 474858
rect 517992 474758 518092 474858
rect 518216 474758 518316 474858
rect 518440 474758 518540 474858
rect 518664 474758 518764 474858
rect 518888 474758 518988 474858
rect 519112 474758 519212 474858
rect 519336 474758 519436 474858
rect 519560 474758 519660 474858
rect 519784 474758 519884 474858
rect 520008 474758 520108 474858
rect 520232 474758 520332 474858
rect 520456 474758 520556 474858
rect 520680 474758 520780 474858
rect 520904 474758 521004 474858
rect 521128 474758 521228 474858
rect 521352 474758 521452 474858
rect 521576 474758 521676 474858
rect 521800 474758 521900 474858
rect 522024 474758 522124 474858
rect 522248 474758 522348 474858
rect 522472 474758 522572 474858
rect 522696 474758 522796 474858
rect 522920 474758 523020 474858
rect 523144 474758 523244 474858
rect 523368 474758 523468 474858
rect 523592 474758 523692 474858
rect 523816 474758 523916 474858
rect 517320 474534 517420 474634
rect 517544 474534 517644 474634
rect 517768 474534 517868 474634
rect 517992 474534 518092 474634
rect 518216 474534 518316 474634
rect 518440 474534 518540 474634
rect 518664 474534 518764 474634
rect 518888 474534 518988 474634
rect 519112 474534 519212 474634
rect 519336 474534 519436 474634
rect 519560 474534 519660 474634
rect 519784 474534 519884 474634
rect 520008 474534 520108 474634
rect 520232 474534 520332 474634
rect 520456 474534 520556 474634
rect 520680 474534 520780 474634
rect 520904 474534 521004 474634
rect 521128 474534 521228 474634
rect 521352 474534 521452 474634
rect 521576 474534 521676 474634
rect 521800 474534 521900 474634
rect 522024 474534 522124 474634
rect 522248 474534 522348 474634
rect 522472 474534 522572 474634
rect 522696 474534 522796 474634
rect 522920 474534 523020 474634
rect 523144 474534 523244 474634
rect 523368 474534 523468 474634
rect 523592 474534 523692 474634
rect 523816 474534 523916 474634
rect 517320 474310 517420 474410
rect 517544 474310 517644 474410
rect 517768 474310 517868 474410
rect 517992 474310 518092 474410
rect 518216 474310 518316 474410
rect 518440 474310 518540 474410
rect 518664 474310 518764 474410
rect 518888 474310 518988 474410
rect 519112 474310 519212 474410
rect 519336 474310 519436 474410
rect 519560 474310 519660 474410
rect 519784 474310 519884 474410
rect 520008 474310 520108 474410
rect 520232 474310 520332 474410
rect 520456 474310 520556 474410
rect 520680 474310 520780 474410
rect 520904 474310 521004 474410
rect 521128 474310 521228 474410
rect 521352 474310 521452 474410
rect 521576 474310 521676 474410
rect 521800 474310 521900 474410
rect 522024 474310 522124 474410
rect 522248 474310 522348 474410
rect 522472 474310 522572 474410
rect 522696 474310 522796 474410
rect 522920 474310 523020 474410
rect 523144 474310 523244 474410
rect 523368 474310 523468 474410
rect 523592 474310 523692 474410
rect 523816 474310 523916 474410
rect 500398 473956 500498 474056
rect 500622 473956 500722 474056
rect 500846 473956 500946 474056
rect 501070 473956 501170 474056
rect 501294 473956 501394 474056
rect 500398 473732 500498 473832
rect 500622 473732 500722 473832
rect 500846 473732 500946 473832
rect 501070 473732 501170 473832
rect 501294 473732 501394 473832
rect 500398 473508 500498 473608
rect 500622 473508 500722 473608
rect 500846 473508 500946 473608
rect 501070 473508 501170 473608
rect 501294 473508 501394 473608
rect 500398 473284 500498 473384
rect 500622 473284 500722 473384
rect 500846 473284 500946 473384
rect 501070 473284 501170 473384
rect 501294 473284 501394 473384
rect 500398 473060 500498 473160
rect 500622 473060 500722 473160
rect 500846 473060 500946 473160
rect 501070 473060 501170 473160
rect 501294 473060 501394 473160
rect 500398 472836 500498 472936
rect 500622 472836 500722 472936
rect 500846 472836 500946 472936
rect 501070 472836 501170 472936
rect 501294 472836 501394 472936
rect 500398 472612 500498 472712
rect 500622 472612 500722 472712
rect 500846 472612 500946 472712
rect 501070 472612 501170 472712
rect 501294 472612 501394 472712
rect 500398 472388 500498 472488
rect 500622 472388 500722 472488
rect 500846 472388 500946 472488
rect 501070 472388 501170 472488
rect 501294 472388 501394 472488
rect 500398 472164 500498 472264
rect 500622 472164 500722 472264
rect 500846 472164 500946 472264
rect 501070 472164 501170 472264
rect 501294 472164 501394 472264
rect 500398 471940 500498 472040
rect 500622 471940 500722 472040
rect 500846 471940 500946 472040
rect 501070 471940 501170 472040
rect 501294 471940 501394 472040
rect 500398 471716 500498 471816
rect 500622 471716 500722 471816
rect 500846 471716 500946 471816
rect 501070 471716 501170 471816
rect 501294 471716 501394 471816
rect 500398 471492 500498 471592
rect 500622 471492 500722 471592
rect 500846 471492 500946 471592
rect 501070 471492 501170 471592
rect 501294 471492 501394 471592
rect 500398 471268 500498 471368
rect 500622 471268 500722 471368
rect 500846 471268 500946 471368
rect 501070 471268 501170 471368
rect 501294 471268 501394 471368
rect 511648 474212 511712 474276
rect 511776 474212 511840 474276
rect 511904 474212 511968 474276
rect 512032 474212 512096 474276
rect 500398 471044 500498 471144
rect 500622 471044 500722 471144
rect 500846 471044 500946 471144
rect 501070 471044 501170 471144
rect 501294 471044 501394 471144
rect 500398 470820 500498 470920
rect 500622 470820 500722 470920
rect 500846 470820 500946 470920
rect 501070 470820 501170 470920
rect 501294 470820 501394 470920
rect 500398 470596 500498 470696
rect 500622 470596 500722 470696
rect 500846 470596 500946 470696
rect 501070 470596 501170 470696
rect 501294 470596 501394 470696
rect 500398 470372 500498 470472
rect 500622 470372 500722 470472
rect 500846 470372 500946 470472
rect 501070 470372 501170 470472
rect 501294 470372 501394 470472
rect 500398 470148 500498 470248
rect 500622 470148 500722 470248
rect 500846 470148 500946 470248
rect 501070 470148 501170 470248
rect 501294 470148 501394 470248
rect 500398 469924 500498 470024
rect 500622 469924 500722 470024
rect 500846 469924 500946 470024
rect 501070 469924 501170 470024
rect 501294 469924 501394 470024
rect 500398 469700 500498 469800
rect 500622 469700 500722 469800
rect 500846 469700 500946 469800
rect 501070 469700 501170 469800
rect 501294 469700 501394 469800
rect 500398 469476 500498 469576
rect 500622 469476 500722 469576
rect 500846 469476 500946 469576
rect 501070 469476 501170 469576
rect 501294 469476 501394 469576
rect 500398 469252 500498 469352
rect 500622 469252 500722 469352
rect 500846 469252 500946 469352
rect 501070 469252 501170 469352
rect 501294 469252 501394 469352
rect 500398 469028 500498 469128
rect 500622 469028 500722 469128
rect 500846 469028 500946 469128
rect 501070 469028 501170 469128
rect 501294 469028 501394 469128
rect 500398 468804 500498 468904
rect 500622 468804 500722 468904
rect 500846 468804 500946 468904
rect 501070 468804 501170 468904
rect 501294 468804 501394 468904
rect 500398 468580 500498 468680
rect 500622 468580 500722 468680
rect 500846 468580 500946 468680
rect 501070 468580 501170 468680
rect 501294 468580 501394 468680
rect 500398 468356 500498 468456
rect 500622 468356 500722 468456
rect 500846 468356 500946 468456
rect 501070 468356 501170 468456
rect 501294 468356 501394 468456
rect 491256 463452 497000 468236
rect 500398 468132 500498 468232
rect 500622 468132 500722 468232
rect 500846 468132 500946 468232
rect 501070 468132 501170 468232
rect 501294 468132 501394 468232
rect 500398 467908 500498 468008
rect 500622 467908 500722 468008
rect 500846 467908 500946 468008
rect 501070 467908 501170 468008
rect 501294 467908 501394 468008
rect 500398 467684 500498 467784
rect 500622 467684 500722 467784
rect 500846 467684 500946 467784
rect 501070 467684 501170 467784
rect 501294 467684 501394 467784
rect 500398 463710 500498 463810
rect 500622 463710 500722 463810
rect 500846 463710 500946 463810
rect 501070 463710 501170 463810
rect 501294 463710 501394 463810
rect 500398 463486 500498 463586
rect 500622 463486 500722 463586
rect 500846 463486 500946 463586
rect 501070 463486 501170 463586
rect 501294 463486 501394 463586
rect 500398 463262 500498 463362
rect 500622 463262 500722 463362
rect 500846 463262 500946 463362
rect 501070 463262 501170 463362
rect 501294 463262 501394 463362
rect 500398 463038 500498 463138
rect 500622 463038 500722 463138
rect 500846 463038 500946 463138
rect 501070 463038 501170 463138
rect 501294 463038 501394 463138
rect 500398 462814 500498 462914
rect 500622 462814 500722 462914
rect 500846 462814 500946 462914
rect 501070 462814 501170 462914
rect 501294 462814 501394 462914
rect 500398 462590 500498 462690
rect 500622 462590 500722 462690
rect 500846 462590 500946 462690
rect 501070 462590 501170 462690
rect 501294 462590 501394 462690
rect 500398 462366 500498 462466
rect 500622 462366 500722 462466
rect 500846 462366 500946 462466
rect 501070 462366 501170 462466
rect 501294 462366 501394 462466
rect 491256 457452 497000 462236
rect 500398 462142 500498 462242
rect 500622 462142 500722 462242
rect 500846 462142 500946 462242
rect 501070 462142 501170 462242
rect 501294 462142 501394 462242
rect 500398 461918 500498 462018
rect 500622 461918 500722 462018
rect 500846 461918 500946 462018
rect 501070 461918 501170 462018
rect 501294 461918 501394 462018
rect 500398 461694 500498 461794
rect 500622 461694 500722 461794
rect 500846 461694 500946 461794
rect 501070 461694 501170 461794
rect 501294 461694 501394 461794
rect 500398 461470 500498 461570
rect 500622 461470 500722 461570
rect 500846 461470 500946 461570
rect 501070 461470 501170 461570
rect 501294 461470 501394 461570
rect 500398 461246 500498 461346
rect 500622 461246 500722 461346
rect 500846 461246 500946 461346
rect 501070 461246 501170 461346
rect 501294 461246 501394 461346
rect 500398 461022 500498 461122
rect 500622 461022 500722 461122
rect 500846 461022 500946 461122
rect 501070 461022 501170 461122
rect 501294 461022 501394 461122
rect 500398 460798 500498 460898
rect 500622 460798 500722 460898
rect 500846 460798 500946 460898
rect 501070 460798 501170 460898
rect 501294 460798 501394 460898
rect 500398 460574 500498 460674
rect 500622 460574 500722 460674
rect 500846 460574 500946 460674
rect 501070 460574 501170 460674
rect 501294 460574 501394 460674
rect 500398 460350 500498 460450
rect 500622 460350 500722 460450
rect 500846 460350 500946 460450
rect 501070 460350 501170 460450
rect 501294 460350 501394 460450
rect 500398 460126 500498 460226
rect 500622 460126 500722 460226
rect 500846 460126 500946 460226
rect 501070 460126 501170 460226
rect 501294 460126 501394 460226
rect 500398 459902 500498 460002
rect 500622 459902 500722 460002
rect 500846 459902 500946 460002
rect 501070 459902 501170 460002
rect 501294 459902 501394 460002
rect 500398 459678 500498 459778
rect 500622 459678 500722 459778
rect 500846 459678 500946 459778
rect 501070 459678 501170 459778
rect 501294 459678 501394 459778
rect 500398 459454 500498 459554
rect 500622 459454 500722 459554
rect 500846 459454 500946 459554
rect 501070 459454 501170 459554
rect 501294 459454 501394 459554
rect 500398 459230 500498 459330
rect 500622 459230 500722 459330
rect 500846 459230 500946 459330
rect 501070 459230 501170 459330
rect 501294 459230 501394 459330
rect 500398 459006 500498 459106
rect 500622 459006 500722 459106
rect 500846 459006 500946 459106
rect 501070 459006 501170 459106
rect 501294 459006 501394 459106
rect 500398 458782 500498 458882
rect 500622 458782 500722 458882
rect 500846 458782 500946 458882
rect 501070 458782 501170 458882
rect 501294 458782 501394 458882
rect 500398 458558 500498 458658
rect 500622 458558 500722 458658
rect 500846 458558 500946 458658
rect 501070 458558 501170 458658
rect 501294 458558 501394 458658
rect 500398 458334 500498 458434
rect 500622 458334 500722 458434
rect 500846 458334 500946 458434
rect 501070 458334 501170 458434
rect 501294 458334 501394 458434
rect 500398 458110 500498 458210
rect 500622 458110 500722 458210
rect 500846 458110 500946 458210
rect 501070 458110 501170 458210
rect 501294 458110 501394 458210
rect 500398 457886 500498 457986
rect 500622 457886 500722 457986
rect 500846 457886 500946 457986
rect 501070 457886 501170 457986
rect 501294 457886 501394 457986
rect 500398 457662 500498 457762
rect 500622 457662 500722 457762
rect 500846 457662 500946 457762
rect 501070 457662 501170 457762
rect 501294 457662 501394 457762
rect 500398 457438 500498 457538
rect 500622 457438 500722 457538
rect 500846 457438 500946 457538
rect 501070 457438 501170 457538
rect 501294 457438 501394 457538
rect 500398 457214 500498 457314
rect 500622 457214 500722 457314
rect 500846 457214 500946 457314
rect 501070 457214 501170 457314
rect 501294 457214 501394 457314
rect 527618 474180 527718 474280
rect 527842 474180 527942 474280
rect 528066 474180 528166 474280
rect 528290 474180 528390 474280
rect 528514 474180 528614 474280
rect 527618 473956 527718 474056
rect 527842 473956 527942 474056
rect 528066 473956 528166 474056
rect 528290 473956 528390 474056
rect 528514 473956 528614 474056
rect 527618 473732 527718 473832
rect 527842 473732 527942 473832
rect 528066 473732 528166 473832
rect 528290 473732 528390 473832
rect 528514 473732 528614 473832
rect 527618 473508 527718 473608
rect 527842 473508 527942 473608
rect 528066 473508 528166 473608
rect 528290 473508 528390 473608
rect 528514 473508 528614 473608
rect 527618 473284 527718 473384
rect 527842 473284 527942 473384
rect 528066 473284 528166 473384
rect 528290 473284 528390 473384
rect 528514 473284 528614 473384
rect 527618 473060 527718 473160
rect 527842 473060 527942 473160
rect 528066 473060 528166 473160
rect 528290 473060 528390 473160
rect 528514 473060 528614 473160
rect 527618 472836 527718 472936
rect 527842 472836 527942 472936
rect 528066 472836 528166 472936
rect 528290 472836 528390 472936
rect 528514 472836 528614 472936
rect 527618 472612 527718 472712
rect 527842 472612 527942 472712
rect 528066 472612 528166 472712
rect 528290 472612 528390 472712
rect 528514 472612 528614 472712
rect 505789 469552 506069 469566
rect 505789 468952 505803 469552
rect 505803 468952 506055 469552
rect 506055 468952 506069 469552
rect 505789 468938 506069 468952
rect 511220 468161 511764 468225
rect 511920 468161 512464 468225
rect 512620 468161 513164 468225
rect 513320 468161 513864 468225
rect 514020 468161 514564 468225
rect 514720 468161 515264 468225
rect 515420 468161 515964 468225
rect 516120 468161 516664 468225
rect 516820 468161 517364 468225
rect 517520 468161 518064 468225
rect 511220 467442 511764 467506
rect 511920 467442 512464 467506
rect 512620 467442 513164 467506
rect 513320 467442 513864 467506
rect 514020 467442 514564 467506
rect 514720 467442 515264 467506
rect 515420 467442 515964 467506
rect 516120 467442 516664 467506
rect 516820 467442 517364 467506
rect 517520 467442 518064 467506
rect 511220 466723 511764 466787
rect 511920 466723 512464 466787
rect 512620 466723 513164 466787
rect 513320 466723 513864 466787
rect 514020 466723 514564 466787
rect 514720 466723 515264 466787
rect 515420 466723 515964 466787
rect 516120 466723 516664 466787
rect 516820 466723 517364 466787
rect 517520 466723 518064 466787
rect 511220 466004 511764 466068
rect 511920 466004 512464 466068
rect 512620 466004 513164 466068
rect 513320 466004 513864 466068
rect 514020 466004 514564 466068
rect 514720 466004 515264 466068
rect 515420 466004 515964 466068
rect 516120 466004 516664 466068
rect 516820 466004 517364 466068
rect 517520 466004 518064 466068
rect 511220 465285 511764 465349
rect 511920 465285 512464 465349
rect 512620 465285 513164 465349
rect 513320 465285 513864 465349
rect 514020 465285 514564 465349
rect 514720 465285 515264 465349
rect 515420 465285 515964 465349
rect 516120 465285 516664 465349
rect 516820 465285 517364 465349
rect 517520 465285 518064 465349
rect 511220 464566 511764 464630
rect 511920 464566 512464 464630
rect 512620 464566 513164 464630
rect 513320 464566 513864 464630
rect 514020 464566 514564 464630
rect 514720 464566 515264 464630
rect 515420 464566 515964 464630
rect 516120 464566 516664 464630
rect 516820 464566 517364 464630
rect 517520 464566 518064 464630
rect 511220 463847 511764 463911
rect 511920 463847 512464 463911
rect 512620 463847 513164 463911
rect 513320 463847 513864 463911
rect 514020 463847 514564 463911
rect 514720 463847 515264 463911
rect 515420 463847 515964 463911
rect 516120 463847 516664 463911
rect 516820 463847 517364 463911
rect 517520 463847 518064 463911
rect 511220 463128 511764 463192
rect 511920 463128 512464 463192
rect 512620 463128 513164 463192
rect 513320 463128 513864 463192
rect 514020 463128 514564 463192
rect 514720 463128 515264 463192
rect 515420 463128 515964 463192
rect 516120 463128 516664 463192
rect 516820 463128 517364 463192
rect 517520 463128 518064 463192
rect 511220 462409 511764 462473
rect 511920 462409 512464 462473
rect 512620 462409 513164 462473
rect 513320 462409 513864 462473
rect 514020 462409 514564 462473
rect 514720 462409 515264 462473
rect 515420 462409 515964 462473
rect 516120 462409 516664 462473
rect 516820 462409 517364 462473
rect 517520 462409 518064 462473
rect 511220 461690 511764 461754
rect 511920 461690 512464 461754
rect 512620 461690 513164 461754
rect 513320 461690 513864 461754
rect 514020 461690 514564 461754
rect 514720 461690 515264 461754
rect 515420 461690 515964 461754
rect 516120 461690 516664 461754
rect 516820 461690 517364 461754
rect 517520 461690 518064 461754
rect 525651 472504 526507 472513
rect 525651 461248 525660 472504
rect 525660 461248 526498 472504
rect 526498 461248 526507 472504
rect 525651 461239 526507 461248
rect 527618 472388 527718 472488
rect 527842 472388 527942 472488
rect 528066 472388 528166 472488
rect 528290 472388 528390 472488
rect 528514 472388 528614 472488
rect 527618 472164 527718 472264
rect 527842 472164 527942 472264
rect 528066 472164 528166 472264
rect 528290 472164 528390 472264
rect 528514 472164 528614 472264
rect 527618 471940 527718 472040
rect 527842 471940 527942 472040
rect 528066 471940 528166 472040
rect 528290 471940 528390 472040
rect 528514 471940 528614 472040
rect 527618 471716 527718 471816
rect 527842 471716 527942 471816
rect 528066 471716 528166 471816
rect 528290 471716 528390 471816
rect 528514 471716 528614 471816
rect 527618 471492 527718 471592
rect 527842 471492 527942 471592
rect 528066 471492 528166 471592
rect 528290 471492 528390 471592
rect 528514 471492 528614 471592
rect 527618 471268 527718 471368
rect 527842 471268 527942 471368
rect 528066 471268 528166 471368
rect 528290 471268 528390 471368
rect 528514 471268 528614 471368
rect 527618 471044 527718 471144
rect 527842 471044 527942 471144
rect 528066 471044 528166 471144
rect 528290 471044 528390 471144
rect 528514 471044 528614 471144
rect 527618 470820 527718 470920
rect 527842 470820 527942 470920
rect 528066 470820 528166 470920
rect 528290 470820 528390 470920
rect 528514 470820 528614 470920
rect 527618 470596 527718 470696
rect 527842 470596 527942 470696
rect 528066 470596 528166 470696
rect 528290 470596 528390 470696
rect 528514 470596 528614 470696
rect 527618 470372 527718 470472
rect 527842 470372 527942 470472
rect 528066 470372 528166 470472
rect 528290 470372 528390 470472
rect 528514 470372 528614 470472
rect 527618 470148 527718 470248
rect 527842 470148 527942 470248
rect 528066 470148 528166 470248
rect 528290 470148 528390 470248
rect 528514 470148 528614 470248
rect 527618 469924 527718 470024
rect 527842 469924 527942 470024
rect 528066 469924 528166 470024
rect 528290 469924 528390 470024
rect 528514 469924 528614 470024
rect 527618 469700 527718 469800
rect 527842 469700 527942 469800
rect 528066 469700 528166 469800
rect 528290 469700 528390 469800
rect 528514 469700 528614 469800
rect 527618 469476 527718 469576
rect 527842 469476 527942 469576
rect 528066 469476 528166 469576
rect 528290 469476 528390 469576
rect 528514 469476 528614 469576
rect 530760 469452 536504 474236
rect 527618 469252 527718 469352
rect 527842 469252 527942 469352
rect 528066 469252 528166 469352
rect 528290 469252 528390 469352
rect 528514 469252 528614 469352
rect 527618 469028 527718 469128
rect 527842 469028 527942 469128
rect 528066 469028 528166 469128
rect 528290 469028 528390 469128
rect 528514 469028 528614 469128
rect 527618 468804 527718 468904
rect 527842 468804 527942 468904
rect 528066 468804 528166 468904
rect 528290 468804 528390 468904
rect 528514 468804 528614 468904
rect 527618 468580 527718 468680
rect 527842 468580 527942 468680
rect 528066 468580 528166 468680
rect 528290 468580 528390 468680
rect 528514 468580 528614 468680
rect 527618 468356 527718 468456
rect 527842 468356 527942 468456
rect 528066 468356 528166 468456
rect 528290 468356 528390 468456
rect 528514 468356 528614 468456
rect 527618 468132 527718 468232
rect 527842 468132 527942 468232
rect 528066 468132 528166 468232
rect 528290 468132 528390 468232
rect 528514 468132 528614 468232
rect 527618 467908 527718 468008
rect 527842 467908 527942 468008
rect 528066 467908 528166 468008
rect 528290 467908 528390 468008
rect 528514 467908 528614 468008
rect 527618 467684 527718 467784
rect 527842 467684 527942 467784
rect 528066 467684 528166 467784
rect 528290 467684 528390 467784
rect 528514 467684 528614 467784
rect 527618 463710 527718 463810
rect 527842 463710 527942 463810
rect 528066 463710 528166 463810
rect 528290 463710 528390 463810
rect 528514 463710 528614 463810
rect 527618 463486 527718 463586
rect 527842 463486 527942 463586
rect 528066 463486 528166 463586
rect 528290 463486 528390 463586
rect 528514 463486 528614 463586
rect 530760 463452 536504 468236
rect 527618 463262 527718 463362
rect 527842 463262 527942 463362
rect 528066 463262 528166 463362
rect 528290 463262 528390 463362
rect 528514 463262 528614 463362
rect 527618 463038 527718 463138
rect 527842 463038 527942 463138
rect 528066 463038 528166 463138
rect 528290 463038 528390 463138
rect 528514 463038 528614 463138
rect 527618 462814 527718 462914
rect 527842 462814 527942 462914
rect 528066 462814 528166 462914
rect 528290 462814 528390 462914
rect 528514 462814 528614 462914
rect 527618 462590 527718 462690
rect 527842 462590 527942 462690
rect 528066 462590 528166 462690
rect 528290 462590 528390 462690
rect 528514 462590 528614 462690
rect 527618 462366 527718 462466
rect 527842 462366 527942 462466
rect 528066 462366 528166 462466
rect 528290 462366 528390 462466
rect 528514 462366 528614 462466
rect 527618 462142 527718 462242
rect 527842 462142 527942 462242
rect 528066 462142 528166 462242
rect 528290 462142 528390 462242
rect 528514 462142 528614 462242
rect 527618 461918 527718 462018
rect 527842 461918 527942 462018
rect 528066 461918 528166 462018
rect 528290 461918 528390 462018
rect 528514 461918 528614 462018
rect 527618 461694 527718 461794
rect 527842 461694 527942 461794
rect 528066 461694 528166 461794
rect 528290 461694 528390 461794
rect 528514 461694 528614 461794
rect 527618 461470 527718 461570
rect 527842 461470 527942 461570
rect 528066 461470 528166 461570
rect 528290 461470 528390 461570
rect 528514 461470 528614 461570
rect 527618 461246 527718 461346
rect 527842 461246 527942 461346
rect 528066 461246 528166 461346
rect 528290 461246 528390 461346
rect 528514 461246 528614 461346
rect 477500 450892 483244 455676
rect 477500 442892 483244 447676
rect 505789 461061 506069 461075
rect 505789 460461 505803 461061
rect 505803 460461 506055 461061
rect 506055 460461 506069 461061
rect 505789 460447 506069 460461
rect 527618 461022 527718 461122
rect 527842 461022 527942 461122
rect 528066 461022 528166 461122
rect 528290 461022 528390 461122
rect 528514 461022 528614 461122
rect 527618 460798 527718 460898
rect 527842 460798 527942 460898
rect 528066 460798 528166 460898
rect 528290 460798 528390 460898
rect 528514 460798 528614 460898
rect 527618 460574 527718 460674
rect 527842 460574 527942 460674
rect 528066 460574 528166 460674
rect 528290 460574 528390 460674
rect 528514 460574 528614 460674
rect 527618 460350 527718 460450
rect 527842 460350 527942 460450
rect 528066 460350 528166 460450
rect 528290 460350 528390 460450
rect 528514 460350 528614 460450
rect 512234 439888 513206 460198
rect 527618 460126 527718 460226
rect 527842 460126 527942 460226
rect 528066 460126 528166 460226
rect 528290 460126 528390 460226
rect 528514 460126 528614 460226
rect 527618 459902 527718 460002
rect 527842 459902 527942 460002
rect 528066 459902 528166 460002
rect 528290 459902 528390 460002
rect 528514 459902 528614 460002
rect 527618 459678 527718 459778
rect 527842 459678 527942 459778
rect 528066 459678 528166 459778
rect 528290 459678 528390 459778
rect 528514 459678 528614 459778
rect 527618 459454 527718 459554
rect 527842 459454 527942 459554
rect 528066 459454 528166 459554
rect 528290 459454 528390 459554
rect 528514 459454 528614 459554
rect 527618 459230 527718 459330
rect 527842 459230 527942 459330
rect 528066 459230 528166 459330
rect 528290 459230 528390 459330
rect 528514 459230 528614 459330
rect 527618 459006 527718 459106
rect 527842 459006 527942 459106
rect 528066 459006 528166 459106
rect 528290 459006 528390 459106
rect 528514 459006 528614 459106
rect 527618 458782 527718 458882
rect 527842 458782 527942 458882
rect 528066 458782 528166 458882
rect 528290 458782 528390 458882
rect 528514 458782 528614 458882
rect 527618 458558 527718 458658
rect 527842 458558 527942 458658
rect 528066 458558 528166 458658
rect 528290 458558 528390 458658
rect 528514 458558 528614 458658
rect 527618 458334 527718 458434
rect 527842 458334 527942 458434
rect 528066 458334 528166 458434
rect 528290 458334 528390 458434
rect 528514 458334 528614 458434
rect 527618 458110 527718 458210
rect 527842 458110 527942 458210
rect 528066 458110 528166 458210
rect 528290 458110 528390 458210
rect 528514 458110 528614 458210
rect 527618 457886 527718 457986
rect 527842 457886 527942 457986
rect 528066 457886 528166 457986
rect 528290 457886 528390 457986
rect 528514 457886 528614 457986
rect 527618 457662 527718 457762
rect 527842 457662 527942 457762
rect 528066 457662 528166 457762
rect 528290 457662 528390 457762
rect 528514 457662 528614 457762
rect 527618 457438 527718 457538
rect 527842 457438 527942 457538
rect 528066 457438 528166 457538
rect 528290 457438 528390 457538
rect 528514 457438 528614 457538
rect 530760 457452 536504 462236
rect 527618 457214 527718 457314
rect 527842 457214 527942 457314
rect 528066 457214 528166 457314
rect 528290 457214 528390 457314
rect 528514 457214 528614 457314
rect 562480 455360 562560 455440
rect 562640 455360 562720 455440
rect 562800 455360 562880 455440
rect 562960 455360 563040 455440
rect 563120 455360 563200 455440
rect 563280 455360 563360 455440
rect 563440 455360 563520 455440
rect 563600 455360 563680 455440
rect 563760 455360 563840 455440
rect 563920 455360 564000 455440
rect 564080 455360 564160 455440
rect 564240 455360 564320 455440
rect 564400 455360 564480 455440
rect 564560 455360 564640 455440
rect 564720 455360 564800 455440
rect 564880 455360 564960 455440
rect 565040 455360 565120 455440
rect 565200 455360 565280 455440
rect 565360 455360 565440 455440
rect 565520 455360 565600 455440
rect 565680 455360 565760 455440
rect 565840 455360 565920 455440
rect 566000 455360 566080 455440
rect 566160 455360 566240 455440
rect 566320 455360 566400 455440
rect 566480 455360 566560 455440
rect 566640 455360 566720 455440
rect 566800 455360 566880 455440
rect 566960 455360 567040 455440
rect 567120 455360 567200 455440
rect 567280 455360 567360 455440
rect 562480 455200 562560 455280
rect 562640 455200 562720 455280
rect 562800 455200 562880 455280
rect 562960 455200 563040 455280
rect 563120 455200 563200 455280
rect 563280 455200 563360 455280
rect 563440 455200 563520 455280
rect 563600 455200 563680 455280
rect 563760 455200 563840 455280
rect 563920 455200 564000 455280
rect 564080 455200 564160 455280
rect 564240 455200 564320 455280
rect 564400 455200 564480 455280
rect 564560 455200 564640 455280
rect 564720 455200 564800 455280
rect 564880 455200 564960 455280
rect 565040 455200 565120 455280
rect 565200 455200 565280 455280
rect 565360 455200 565440 455280
rect 565520 455200 565600 455280
rect 565680 455200 565760 455280
rect 565840 455200 565920 455280
rect 566000 455200 566080 455280
rect 566160 455200 566240 455280
rect 566320 455200 566400 455280
rect 566480 455200 566560 455280
rect 566640 455200 566720 455280
rect 566800 455200 566880 455280
rect 566960 455200 567040 455280
rect 567120 455200 567200 455280
rect 567280 455200 567360 455280
rect 572640 455360 572720 455440
rect 572800 455360 572880 455440
rect 572960 455360 573040 455440
rect 573120 455360 573200 455440
rect 573280 455360 573360 455440
rect 573440 455360 573520 455440
rect 573600 455360 573680 455440
rect 573760 455360 573840 455440
rect 573920 455360 574000 455440
rect 574080 455360 574160 455440
rect 574240 455360 574320 455440
rect 574400 455360 574480 455440
rect 574560 455360 574640 455440
rect 574720 455360 574800 455440
rect 574880 455360 574960 455440
rect 575040 455360 575120 455440
rect 575200 455360 575280 455440
rect 575360 455360 575440 455440
rect 575520 455360 575600 455440
rect 575680 455360 575760 455440
rect 575840 455360 575920 455440
rect 576000 455360 576080 455440
rect 576160 455360 576240 455440
rect 576320 455360 576400 455440
rect 576480 455360 576560 455440
rect 576640 455360 576720 455440
rect 576800 455360 576880 455440
rect 576960 455360 577040 455440
rect 577120 455360 577200 455440
rect 577280 455360 577360 455440
rect 577440 455360 577520 455440
rect 572640 455200 572720 455280
rect 572800 455200 572880 455280
rect 572960 455200 573040 455280
rect 573120 455200 573200 455280
rect 573280 455200 573360 455280
rect 573440 455200 573520 455280
rect 573600 455200 573680 455280
rect 573760 455200 573840 455280
rect 573920 455200 574000 455280
rect 574080 455200 574160 455280
rect 574240 455200 574320 455280
rect 574400 455200 574480 455280
rect 574560 455200 574640 455280
rect 574720 455200 574800 455280
rect 574880 455200 574960 455280
rect 575040 455200 575120 455280
rect 575200 455200 575280 455280
rect 575360 455200 575440 455280
rect 575520 455200 575600 455280
rect 575680 455200 575760 455280
rect 575840 455200 575920 455280
rect 576000 455200 576080 455280
rect 576160 455200 576240 455280
rect 576320 455200 576400 455280
rect 576480 455200 576560 455280
rect 576640 455200 576720 455280
rect 576800 455200 576880 455280
rect 576960 455200 577040 455280
rect 577120 455200 577200 455280
rect 577280 455200 577360 455280
rect 577440 455200 577520 455280
rect 513720 453556 513920 453756
rect 514154 453556 514354 453756
rect 514588 453556 514788 453756
rect 513720 453122 513920 453322
rect 514154 453122 514354 453322
rect 514588 453122 514788 453322
rect 513720 452688 513920 452888
rect 514154 452688 514354 452888
rect 514588 452688 514788 452888
rect 513720 452254 513920 452454
rect 514154 452254 514354 452454
rect 514588 452254 514788 452454
rect 513720 451820 513920 452020
rect 514154 451820 514354 452020
rect 514588 451820 514788 452020
rect 513720 451386 513920 451586
rect 514154 451386 514354 451586
rect 514588 451386 514788 451586
rect 513720 450952 513920 451152
rect 514154 450952 514354 451152
rect 514588 450952 514788 451152
rect 513720 450518 513920 450718
rect 514154 450518 514354 450718
rect 514588 450518 514788 450718
rect 513720 450084 513920 450284
rect 514154 450084 514354 450284
rect 514588 450084 514788 450284
rect 513720 449650 513920 449850
rect 514154 449650 514354 449850
rect 514588 449650 514788 449850
rect 513720 449216 513920 449416
rect 514154 449216 514354 449416
rect 514588 449216 514788 449416
rect 514588 448816 514788 449016
rect 514588 448416 514788 448616
rect 514588 448016 514788 448216
rect 514588 447616 514788 447816
rect 514588 447216 514788 447416
rect 514588 446816 514788 447016
rect 514588 446416 514788 446616
rect 514588 446016 514788 446216
rect 514588 445616 514788 445816
rect 514588 444016 514788 444216
rect 514588 443616 514788 443816
rect 514588 443216 514788 443416
rect 514588 442816 514788 443016
rect 514588 442416 514788 442616
rect 514588 442016 514788 442216
rect 514588 441616 514788 441816
rect 514588 441216 514788 441416
rect 514588 440816 514788 441016
rect 500418 437440 500518 437540
rect 500642 437440 500742 437540
rect 500866 437440 500966 437540
rect 501090 437440 501190 437540
rect 501314 437440 501414 437540
rect 500418 437216 500518 437316
rect 500642 437216 500742 437316
rect 500866 437216 500966 437316
rect 501090 437216 501190 437316
rect 501314 437216 501414 437316
rect 500418 436992 500518 437092
rect 500642 436992 500742 437092
rect 500866 436992 500966 437092
rect 501090 436992 501190 437092
rect 501314 436992 501414 437092
rect 500418 436768 500518 436868
rect 500642 436768 500742 436868
rect 500866 436768 500966 436868
rect 501090 436768 501190 436868
rect 501314 436768 501414 436868
rect 491260 431892 497004 436676
rect 500418 436544 500518 436644
rect 500642 436544 500742 436644
rect 500866 436544 500966 436644
rect 501090 436544 501190 436644
rect 501314 436544 501414 436644
rect 500418 436320 500518 436420
rect 500642 436320 500742 436420
rect 500866 436320 500966 436420
rect 501090 436320 501190 436420
rect 501314 436320 501414 436420
rect 500418 436096 500518 436196
rect 500642 436096 500742 436196
rect 500866 436096 500966 436196
rect 501090 436096 501190 436196
rect 501314 436096 501414 436196
rect 500418 435872 500518 435972
rect 500642 435872 500742 435972
rect 500866 435872 500966 435972
rect 501090 435872 501190 435972
rect 501314 435872 501414 435972
rect 500418 435648 500518 435748
rect 500642 435648 500742 435748
rect 500866 435648 500966 435748
rect 501090 435648 501190 435748
rect 501314 435648 501414 435748
rect 500418 435424 500518 435524
rect 500642 435424 500742 435524
rect 500866 435424 500966 435524
rect 501090 435424 501190 435524
rect 501314 435424 501414 435524
rect 500418 435200 500518 435300
rect 500642 435200 500742 435300
rect 500866 435200 500966 435300
rect 501090 435200 501190 435300
rect 501314 435200 501414 435300
rect 500418 434976 500518 435076
rect 500642 434976 500742 435076
rect 500866 434976 500966 435076
rect 501090 434976 501190 435076
rect 501314 434976 501414 435076
rect 500418 434752 500518 434852
rect 500642 434752 500742 434852
rect 500866 434752 500966 434852
rect 501090 434752 501190 434852
rect 501314 434752 501414 434852
rect 500418 434528 500518 434628
rect 500642 434528 500742 434628
rect 500866 434528 500966 434628
rect 501090 434528 501190 434628
rect 501314 434528 501414 434628
rect 500418 434304 500518 434404
rect 500642 434304 500742 434404
rect 500866 434304 500966 434404
rect 501090 434304 501190 434404
rect 501314 434304 501414 434404
rect 500418 434080 500518 434180
rect 500642 434080 500742 434180
rect 500866 434080 500966 434180
rect 501090 434080 501190 434180
rect 501314 434080 501414 434180
rect 500418 433856 500518 433956
rect 500642 433856 500742 433956
rect 500866 433856 500966 433956
rect 501090 433856 501190 433956
rect 501314 433856 501414 433956
rect 500418 433632 500518 433732
rect 500642 433632 500742 433732
rect 500866 433632 500966 433732
rect 501090 433632 501190 433732
rect 501314 433632 501414 433732
rect 500418 433408 500518 433508
rect 500642 433408 500742 433508
rect 500866 433408 500966 433508
rect 501090 433408 501190 433508
rect 501314 433408 501414 433508
rect 500418 433184 500518 433284
rect 500642 433184 500742 433284
rect 500866 433184 500966 433284
rect 501090 433184 501190 433284
rect 501314 433184 501414 433284
rect 500418 432960 500518 433060
rect 500642 432960 500742 433060
rect 500866 432960 500966 433060
rect 501090 432960 501190 433060
rect 501314 432960 501414 433060
rect 500418 432736 500518 432836
rect 500642 432736 500742 432836
rect 500866 432736 500966 432836
rect 501090 432736 501190 432836
rect 501314 432736 501414 432836
rect 500418 432512 500518 432612
rect 500642 432512 500742 432612
rect 500866 432512 500966 432612
rect 501090 432512 501190 432612
rect 501314 432512 501414 432612
rect 500418 432288 500518 432388
rect 500642 432288 500742 432388
rect 500866 432288 500966 432388
rect 501090 432288 501190 432388
rect 501314 432288 501414 432388
rect 500418 432064 500518 432164
rect 500642 432064 500742 432164
rect 500866 432064 500966 432164
rect 501090 432064 501190 432164
rect 501314 432064 501414 432164
rect 500418 431840 500518 431940
rect 500642 431840 500742 431940
rect 500866 431840 500966 431940
rect 501090 431840 501190 431940
rect 501314 431840 501414 431940
rect 500418 431616 500518 431716
rect 500642 431616 500742 431716
rect 500866 431616 500966 431716
rect 501090 431616 501190 431716
rect 501314 431616 501414 431716
rect 500418 431392 500518 431492
rect 500642 431392 500742 431492
rect 500866 431392 500966 431492
rect 501090 431392 501190 431492
rect 501314 431392 501414 431492
rect 500418 431168 500518 431268
rect 500642 431168 500742 431268
rect 500866 431168 500966 431268
rect 501090 431168 501190 431268
rect 501314 431168 501414 431268
rect 527638 437440 527738 437540
rect 527862 437440 527962 437540
rect 528086 437440 528186 437540
rect 528310 437440 528410 437540
rect 528534 437440 528634 437540
rect 527638 437216 527738 437316
rect 527862 437216 527962 437316
rect 528086 437216 528186 437316
rect 528310 437216 528410 437316
rect 528534 437216 528634 437316
rect 527638 436992 527738 437092
rect 527862 436992 527962 437092
rect 528086 436992 528186 437092
rect 528310 436992 528410 437092
rect 528534 436992 528634 437092
rect 527638 436768 527738 436868
rect 527862 436768 527962 436868
rect 528086 436768 528186 436868
rect 528310 436768 528410 436868
rect 528534 436768 528634 436868
rect 527638 436544 527738 436644
rect 527862 436544 527962 436644
rect 528086 436544 528186 436644
rect 528310 436544 528410 436644
rect 528534 436544 528634 436644
rect 527638 436320 527738 436420
rect 527862 436320 527962 436420
rect 528086 436320 528186 436420
rect 528310 436320 528410 436420
rect 528534 436320 528634 436420
rect 527638 436096 527738 436196
rect 527862 436096 527962 436196
rect 528086 436096 528186 436196
rect 528310 436096 528410 436196
rect 528534 436096 528634 436196
rect 527638 435872 527738 435972
rect 527862 435872 527962 435972
rect 528086 435872 528186 435972
rect 528310 435872 528410 435972
rect 528534 435872 528634 435972
rect 527638 435648 527738 435748
rect 527862 435648 527962 435748
rect 528086 435648 528186 435748
rect 528310 435648 528410 435748
rect 528534 435648 528634 435748
rect 527638 435424 527738 435524
rect 527862 435424 527962 435524
rect 528086 435424 528186 435524
rect 528310 435424 528410 435524
rect 528534 435424 528634 435524
rect 527638 435200 527738 435300
rect 527862 435200 527962 435300
rect 528086 435200 528186 435300
rect 528310 435200 528410 435300
rect 528534 435200 528634 435300
rect 527638 434976 527738 435076
rect 527862 434976 527962 435076
rect 528086 434976 528186 435076
rect 528310 434976 528410 435076
rect 528534 434976 528634 435076
rect 527638 434752 527738 434852
rect 527862 434752 527962 434852
rect 528086 434752 528186 434852
rect 528310 434752 528410 434852
rect 528534 434752 528634 434852
rect 527638 434528 527738 434628
rect 527862 434528 527962 434628
rect 528086 434528 528186 434628
rect 528310 434528 528410 434628
rect 528534 434528 528634 434628
rect 527638 434304 527738 434404
rect 527862 434304 527962 434404
rect 528086 434304 528186 434404
rect 528310 434304 528410 434404
rect 528534 434304 528634 434404
rect 527638 434080 527738 434180
rect 527862 434080 527962 434180
rect 528086 434080 528186 434180
rect 528310 434080 528410 434180
rect 528534 434080 528634 434180
rect 527638 433856 527738 433956
rect 527862 433856 527962 433956
rect 528086 433856 528186 433956
rect 528310 433856 528410 433956
rect 528534 433856 528634 433956
rect 527638 433632 527738 433732
rect 527862 433632 527962 433732
rect 528086 433632 528186 433732
rect 528310 433632 528410 433732
rect 528534 433632 528634 433732
rect 527638 433408 527738 433508
rect 527862 433408 527962 433508
rect 528086 433408 528186 433508
rect 528310 433408 528410 433508
rect 528534 433408 528634 433508
rect 527638 433184 527738 433284
rect 527862 433184 527962 433284
rect 528086 433184 528186 433284
rect 528310 433184 528410 433284
rect 528534 433184 528634 433284
rect 527638 432960 527738 433060
rect 527862 432960 527962 433060
rect 528086 432960 528186 433060
rect 528310 432960 528410 433060
rect 528534 432960 528634 433060
rect 527638 432736 527738 432836
rect 527862 432736 527962 432836
rect 528086 432736 528186 432836
rect 528310 432736 528410 432836
rect 528534 432736 528634 432836
rect 527638 432512 527738 432612
rect 527862 432512 527962 432612
rect 528086 432512 528186 432612
rect 528310 432512 528410 432612
rect 528534 432512 528634 432612
rect 527638 432288 527738 432388
rect 527862 432288 527962 432388
rect 528086 432288 528186 432388
rect 528310 432288 528410 432388
rect 528534 432288 528634 432388
rect 527638 432064 527738 432164
rect 527862 432064 527962 432164
rect 528086 432064 528186 432164
rect 528310 432064 528410 432164
rect 528534 432064 528634 432164
rect 527638 431840 527738 431940
rect 527862 431840 527962 431940
rect 528086 431840 528186 431940
rect 528310 431840 528410 431940
rect 528534 431840 528634 431940
rect 531080 431892 536824 436676
rect 527638 431616 527738 431716
rect 527862 431616 527962 431716
rect 528086 431616 528186 431716
rect 528310 431616 528410 431716
rect 528534 431616 528634 431716
rect 527638 431392 527738 431492
rect 527862 431392 527962 431492
rect 528086 431392 528186 431492
rect 528310 431392 528410 431492
rect 528534 431392 528634 431492
rect 527638 431168 527738 431268
rect 527862 431168 527962 431268
rect 528086 431168 528186 431268
rect 528310 431168 528410 431268
rect 528534 431168 528634 431268
rect 500418 430944 500518 431044
rect 500642 430944 500742 431044
rect 500866 430944 500966 431044
rect 501090 430944 501190 431044
rect 501314 430944 501414 431044
rect 503920 430926 504020 431026
rect 504144 430926 504244 431026
rect 504368 430926 504468 431026
rect 504592 430926 504692 431026
rect 504816 430926 504916 431026
rect 505040 430926 505140 431026
rect 505264 430926 505364 431026
rect 505488 430926 505588 431026
rect 505712 430926 505812 431026
rect 505936 430926 506036 431026
rect 506160 430926 506260 431026
rect 506384 430926 506484 431026
rect 506608 430926 506708 431026
rect 506832 430926 506932 431026
rect 507056 430926 507156 431026
rect 507280 430926 507380 431026
rect 507504 430926 507604 431026
rect 507728 430926 507828 431026
rect 507952 430926 508052 431026
rect 508176 430926 508276 431026
rect 508400 430926 508500 431026
rect 508624 430926 508724 431026
rect 508848 430926 508948 431026
rect 509072 430926 509172 431026
rect 509296 430926 509396 431026
rect 509520 430926 509620 431026
rect 509744 430926 509844 431026
rect 509968 430926 510068 431026
rect 510192 430926 510292 431026
rect 510416 430926 510516 431026
rect 503920 430702 504020 430802
rect 504144 430702 504244 430802
rect 504368 430702 504468 430802
rect 504592 430702 504692 430802
rect 504816 430702 504916 430802
rect 505040 430702 505140 430802
rect 505264 430702 505364 430802
rect 505488 430702 505588 430802
rect 505712 430702 505812 430802
rect 505936 430702 506036 430802
rect 506160 430702 506260 430802
rect 506384 430702 506484 430802
rect 506608 430702 506708 430802
rect 506832 430702 506932 430802
rect 507056 430702 507156 430802
rect 507280 430702 507380 430802
rect 507504 430702 507604 430802
rect 507728 430702 507828 430802
rect 507952 430702 508052 430802
rect 508176 430702 508276 430802
rect 508400 430702 508500 430802
rect 508624 430702 508724 430802
rect 508848 430702 508948 430802
rect 509072 430702 509172 430802
rect 509296 430702 509396 430802
rect 509520 430702 509620 430802
rect 509744 430702 509844 430802
rect 509968 430702 510068 430802
rect 510192 430702 510292 430802
rect 510416 430702 510516 430802
rect 503920 430478 504020 430578
rect 504144 430478 504244 430578
rect 504368 430478 504468 430578
rect 504592 430478 504692 430578
rect 504816 430478 504916 430578
rect 505040 430478 505140 430578
rect 505264 430478 505364 430578
rect 505488 430478 505588 430578
rect 505712 430478 505812 430578
rect 505936 430478 506036 430578
rect 506160 430478 506260 430578
rect 506384 430478 506484 430578
rect 506608 430478 506708 430578
rect 506832 430478 506932 430578
rect 507056 430478 507156 430578
rect 507280 430478 507380 430578
rect 507504 430478 507604 430578
rect 507728 430478 507828 430578
rect 507952 430478 508052 430578
rect 508176 430478 508276 430578
rect 508400 430478 508500 430578
rect 508624 430478 508724 430578
rect 508848 430478 508948 430578
rect 509072 430478 509172 430578
rect 509296 430478 509396 430578
rect 509520 430478 509620 430578
rect 509744 430478 509844 430578
rect 509968 430478 510068 430578
rect 510192 430478 510292 430578
rect 510416 430478 510516 430578
rect 503920 430254 504020 430354
rect 504144 430254 504244 430354
rect 504368 430254 504468 430354
rect 504592 430254 504692 430354
rect 504816 430254 504916 430354
rect 505040 430254 505140 430354
rect 505264 430254 505364 430354
rect 505488 430254 505588 430354
rect 505712 430254 505812 430354
rect 505936 430254 506036 430354
rect 506160 430254 506260 430354
rect 506384 430254 506484 430354
rect 506608 430254 506708 430354
rect 506832 430254 506932 430354
rect 507056 430254 507156 430354
rect 507280 430254 507380 430354
rect 507504 430254 507604 430354
rect 507728 430254 507828 430354
rect 507952 430254 508052 430354
rect 508176 430254 508276 430354
rect 508400 430254 508500 430354
rect 508624 430254 508724 430354
rect 508848 430254 508948 430354
rect 509072 430254 509172 430354
rect 509296 430254 509396 430354
rect 509520 430254 509620 430354
rect 509744 430254 509844 430354
rect 509968 430254 510068 430354
rect 510192 430254 510292 430354
rect 510416 430254 510516 430354
rect 503920 430030 504020 430130
rect 504144 430030 504244 430130
rect 504368 430030 504468 430130
rect 504592 430030 504692 430130
rect 504816 430030 504916 430130
rect 505040 430030 505140 430130
rect 505264 430030 505364 430130
rect 505488 430030 505588 430130
rect 505712 430030 505812 430130
rect 505936 430030 506036 430130
rect 506160 430030 506260 430130
rect 506384 430030 506484 430130
rect 506608 430030 506708 430130
rect 506832 430030 506932 430130
rect 507056 430030 507156 430130
rect 507280 430030 507380 430130
rect 507504 430030 507604 430130
rect 507728 430030 507828 430130
rect 507952 430030 508052 430130
rect 508176 430030 508276 430130
rect 508400 430030 508500 430130
rect 508624 430030 508724 430130
rect 508848 430030 508948 430130
rect 509072 430030 509172 430130
rect 509296 430030 509396 430130
rect 509520 430030 509620 430130
rect 509744 430030 509844 430130
rect 509968 430030 510068 430130
rect 510192 430030 510292 430130
rect 510416 430030 510516 430130
rect 517320 430926 517420 431026
rect 517544 430926 517644 431026
rect 517768 430926 517868 431026
rect 517992 430926 518092 431026
rect 518216 430926 518316 431026
rect 518440 430926 518540 431026
rect 518664 430926 518764 431026
rect 518888 430926 518988 431026
rect 519112 430926 519212 431026
rect 519336 430926 519436 431026
rect 519560 430926 519660 431026
rect 519784 430926 519884 431026
rect 520008 430926 520108 431026
rect 520232 430926 520332 431026
rect 520456 430926 520556 431026
rect 520680 430926 520780 431026
rect 520904 430926 521004 431026
rect 521128 430926 521228 431026
rect 521352 430926 521452 431026
rect 521576 430926 521676 431026
rect 521800 430926 521900 431026
rect 522024 430926 522124 431026
rect 522248 430926 522348 431026
rect 522472 430926 522572 431026
rect 522696 430926 522796 431026
rect 522920 430926 523020 431026
rect 523144 430926 523244 431026
rect 523368 430926 523468 431026
rect 523592 430926 523692 431026
rect 523816 430926 523916 431026
rect 517320 430702 517420 430802
rect 517544 430702 517644 430802
rect 517768 430702 517868 430802
rect 517992 430702 518092 430802
rect 518216 430702 518316 430802
rect 518440 430702 518540 430802
rect 518664 430702 518764 430802
rect 518888 430702 518988 430802
rect 519112 430702 519212 430802
rect 519336 430702 519436 430802
rect 519560 430702 519660 430802
rect 519784 430702 519884 430802
rect 520008 430702 520108 430802
rect 520232 430702 520332 430802
rect 520456 430702 520556 430802
rect 520680 430702 520780 430802
rect 520904 430702 521004 430802
rect 521128 430702 521228 430802
rect 521352 430702 521452 430802
rect 521576 430702 521676 430802
rect 521800 430702 521900 430802
rect 522024 430702 522124 430802
rect 522248 430702 522348 430802
rect 522472 430702 522572 430802
rect 522696 430702 522796 430802
rect 522920 430702 523020 430802
rect 523144 430702 523244 430802
rect 523368 430702 523468 430802
rect 523592 430702 523692 430802
rect 523816 430702 523916 430802
rect 527638 430944 527738 431044
rect 527862 430944 527962 431044
rect 528086 430944 528186 431044
rect 528310 430944 528410 431044
rect 528534 430944 528634 431044
rect 517320 430478 517420 430578
rect 517544 430478 517644 430578
rect 517768 430478 517868 430578
rect 517992 430478 518092 430578
rect 518216 430478 518316 430578
rect 518440 430478 518540 430578
rect 518664 430478 518764 430578
rect 518888 430478 518988 430578
rect 519112 430478 519212 430578
rect 519336 430478 519436 430578
rect 519560 430478 519660 430578
rect 519784 430478 519884 430578
rect 520008 430478 520108 430578
rect 520232 430478 520332 430578
rect 520456 430478 520556 430578
rect 520680 430478 520780 430578
rect 520904 430478 521004 430578
rect 521128 430478 521228 430578
rect 521352 430478 521452 430578
rect 521576 430478 521676 430578
rect 521800 430478 521900 430578
rect 522024 430478 522124 430578
rect 522248 430478 522348 430578
rect 522472 430478 522572 430578
rect 522696 430478 522796 430578
rect 522920 430478 523020 430578
rect 523144 430478 523244 430578
rect 523368 430478 523468 430578
rect 523592 430478 523692 430578
rect 523816 430478 523916 430578
rect 517320 430254 517420 430354
rect 517544 430254 517644 430354
rect 517768 430254 517868 430354
rect 517992 430254 518092 430354
rect 518216 430254 518316 430354
rect 518440 430254 518540 430354
rect 518664 430254 518764 430354
rect 518888 430254 518988 430354
rect 519112 430254 519212 430354
rect 519336 430254 519436 430354
rect 519560 430254 519660 430354
rect 519784 430254 519884 430354
rect 520008 430254 520108 430354
rect 520232 430254 520332 430354
rect 520456 430254 520556 430354
rect 520680 430254 520780 430354
rect 520904 430254 521004 430354
rect 521128 430254 521228 430354
rect 521352 430254 521452 430354
rect 521576 430254 521676 430354
rect 521800 430254 521900 430354
rect 522024 430254 522124 430354
rect 522248 430254 522348 430354
rect 522472 430254 522572 430354
rect 522696 430254 522796 430354
rect 522920 430254 523020 430354
rect 523144 430254 523244 430354
rect 523368 430254 523468 430354
rect 523592 430254 523692 430354
rect 523816 430254 523916 430354
rect 517320 430030 517420 430130
rect 517544 430030 517644 430130
rect 517768 430030 517868 430130
rect 517992 430030 518092 430130
rect 518216 430030 518316 430130
rect 518440 430030 518540 430130
rect 518664 430030 518764 430130
rect 518888 430030 518988 430130
rect 519112 430030 519212 430130
rect 519336 430030 519436 430130
rect 519560 430030 519660 430130
rect 519784 430030 519884 430130
rect 520008 430030 520108 430130
rect 520232 430030 520332 430130
rect 520456 430030 520556 430130
rect 520680 430030 520780 430130
rect 520904 430030 521004 430130
rect 521128 430030 521228 430130
rect 521352 430030 521452 430130
rect 521576 430030 521676 430130
rect 521800 430030 521900 430130
rect 522024 430030 522124 430130
rect 522248 430030 522348 430130
rect 522472 430030 522572 430130
rect 522696 430030 522796 430130
rect 522920 430030 523020 430130
rect 523144 430030 523244 430130
rect 523368 430030 523468 430130
rect 523592 430030 523692 430130
rect 523816 430030 523916 430130
rect 572772 426216 573008 426452
rect 573244 426216 573480 426452
rect 573716 426216 573952 426452
rect 574188 426216 574424 426452
rect 574660 426216 574896 426452
rect 575132 426216 575368 426452
rect 575604 426216 575840 426452
rect 576076 426216 576312 426452
rect 576548 426216 576784 426452
rect 577020 426216 577256 426452
rect 491138 421216 496882 426000
rect 504338 421216 510082 426000
rect 517738 421216 523482 426000
rect 531138 421216 536882 426000
rect 572772 425744 573008 425980
rect 573244 425744 573480 425980
rect 573716 425744 573952 425980
rect 574188 425744 574424 425980
rect 574660 425744 574896 425980
rect 575132 425744 575368 425980
rect 575604 425744 575840 425980
rect 576076 425744 576312 425980
rect 576548 425744 576784 425980
rect 577020 425744 577256 425980
rect 572772 425272 573008 425508
rect 573244 425272 573480 425508
rect 573716 425272 573952 425508
rect 574188 425272 574424 425508
rect 574660 425272 574896 425508
rect 575132 425272 575368 425508
rect 575604 425272 575840 425508
rect 576076 425272 576312 425508
rect 576548 425272 576784 425508
rect 577020 425272 577256 425508
rect 572772 424800 573008 425036
rect 573244 424800 573480 425036
rect 573716 424800 573952 425036
rect 574188 424800 574424 425036
rect 574660 424800 574896 425036
rect 575132 424800 575368 425036
rect 575604 424800 575840 425036
rect 576076 424800 576312 425036
rect 576548 424800 576784 425036
rect 577020 424800 577256 425036
rect 572772 424328 573008 424564
rect 573244 424328 573480 424564
rect 573716 424328 573952 424564
rect 574188 424328 574424 424564
rect 574660 424328 574896 424564
rect 575132 424328 575368 424564
rect 575604 424328 575840 424564
rect 576076 424328 576312 424564
rect 576548 424328 576784 424564
rect 577020 424328 577256 424564
rect 572772 423856 573008 424092
rect 573244 423856 573480 424092
rect 573716 423856 573952 424092
rect 574188 423856 574424 424092
rect 574660 423856 574896 424092
rect 575132 423856 575368 424092
rect 575604 423856 575840 424092
rect 576076 423856 576312 424092
rect 576548 423856 576784 424092
rect 577020 423856 577256 424092
rect 572772 423384 573008 423620
rect 573244 423384 573480 423620
rect 573716 423384 573952 423620
rect 574188 423384 574424 423620
rect 574660 423384 574896 423620
rect 575132 423384 575368 423620
rect 575604 423384 575840 423620
rect 576076 423384 576312 423620
rect 576548 423384 576784 423620
rect 577020 423384 577256 423620
rect 572772 422912 573008 423148
rect 573244 422912 573480 423148
rect 573716 422912 573952 423148
rect 574188 422912 574424 423148
rect 574660 422912 574896 423148
rect 575132 422912 575368 423148
rect 575604 422912 575840 423148
rect 576076 422912 576312 423148
rect 576548 422912 576784 423148
rect 577020 422912 577256 423148
rect 572772 422440 573008 422676
rect 573244 422440 573480 422676
rect 573716 422440 573952 422676
rect 574188 422440 574424 422676
rect 574660 422440 574896 422676
rect 575132 422440 575368 422676
rect 575604 422440 575840 422676
rect 576076 422440 576312 422676
rect 576548 422440 576784 422676
rect 577020 422440 577256 422676
rect 572772 421968 573008 422204
rect 573244 421968 573480 422204
rect 573716 421968 573952 422204
rect 574188 421968 574424 422204
rect 574660 421968 574896 422204
rect 575132 421968 575368 422204
rect 575604 421968 575840 422204
rect 576076 421968 576312 422204
rect 576548 421968 576784 422204
rect 577020 421968 577256 422204
rect 572772 421496 573008 421732
rect 573244 421496 573480 421732
rect 573716 421496 573952 421732
rect 574188 421496 574424 421732
rect 574660 421496 574896 421732
rect 575132 421496 575368 421732
rect 575604 421496 575840 421732
rect 576076 421496 576312 421732
rect 576548 421496 576784 421732
rect 577020 421496 577256 421732
rect 572772 421024 573008 421260
rect 573244 421024 573480 421260
rect 573716 421024 573952 421260
rect 574188 421024 574424 421260
rect 574660 421024 574896 421260
rect 575132 421024 575368 421260
rect 575604 421024 575840 421260
rect 576076 421024 576312 421260
rect 576548 421024 576784 421260
rect 577020 421024 577256 421260
rect 572772 420552 573008 420788
rect 573244 420552 573480 420788
rect 573716 420552 573952 420788
rect 574188 420552 574424 420788
rect 574660 420552 574896 420788
rect 575132 420552 575368 420788
rect 575604 420552 575840 420788
rect 576076 420552 576312 420788
rect 576548 420552 576784 420788
rect 577020 420552 577256 420788
rect 477192 377600 477428 377836
rect 477664 377600 477900 377836
rect 478136 377600 478372 377836
rect 478608 377600 478844 377836
rect 479080 377600 479316 377836
rect 479552 377600 479788 377836
rect 480024 377600 480260 377836
rect 480496 377600 480732 377836
rect 480968 377600 481204 377836
rect 481440 377600 481676 377836
rect 481912 377600 482148 377836
rect 482384 377600 482620 377836
rect 482856 377600 483092 377836
rect 483328 377600 483564 377836
rect 562624 377364 562860 377600
rect 563096 377364 563332 377600
rect 563568 377364 563804 377600
rect 564040 377364 564276 377600
rect 564512 377364 564748 377600
rect 564984 377364 565220 377600
rect 565456 377364 565692 377600
rect 565928 377364 566164 377600
rect 566400 377364 566636 377600
rect 566872 377364 567108 377600
rect 477192 377128 477428 377364
rect 477664 377128 477900 377364
rect 478136 377128 478372 377364
rect 478608 377128 478844 377364
rect 479080 377128 479316 377364
rect 479552 377128 479788 377364
rect 480024 377128 480260 377364
rect 480496 377128 480732 377364
rect 480968 377128 481204 377364
rect 481440 377128 481676 377364
rect 481912 377128 482148 377364
rect 482384 377128 482620 377364
rect 482856 377128 483092 377364
rect 483328 377128 483564 377364
rect 562624 376892 562860 377128
rect 563096 376892 563332 377128
rect 563568 376892 563804 377128
rect 564040 376892 564276 377128
rect 564512 376892 564748 377128
rect 564984 376892 565220 377128
rect 565456 376892 565692 377128
rect 565928 376892 566164 377128
rect 566400 376892 566636 377128
rect 566872 376892 567108 377128
rect 477192 376656 477428 376892
rect 477664 376656 477900 376892
rect 478136 376656 478372 376892
rect 478608 376656 478844 376892
rect 479080 376656 479316 376892
rect 479552 376656 479788 376892
rect 480024 376656 480260 376892
rect 480496 376656 480732 376892
rect 480968 376656 481204 376892
rect 481440 376656 481676 376892
rect 481912 376656 482148 376892
rect 482384 376656 482620 376892
rect 482856 376656 483092 376892
rect 483328 376656 483564 376892
rect 562624 376420 562860 376656
rect 563096 376420 563332 376656
rect 563568 376420 563804 376656
rect 564040 376420 564276 376656
rect 564512 376420 564748 376656
rect 564984 376420 565220 376656
rect 565456 376420 565692 376656
rect 565928 376420 566164 376656
rect 566400 376420 566636 376656
rect 566872 376420 567108 376656
rect 477192 376184 477428 376420
rect 477664 376184 477900 376420
rect 478136 376184 478372 376420
rect 478608 376184 478844 376420
rect 479080 376184 479316 376420
rect 479552 376184 479788 376420
rect 480024 376184 480260 376420
rect 480496 376184 480732 376420
rect 480968 376184 481204 376420
rect 481440 376184 481676 376420
rect 481912 376184 482148 376420
rect 482384 376184 482620 376420
rect 482856 376184 483092 376420
rect 483328 376184 483564 376420
rect 562624 375948 562860 376184
rect 563096 375948 563332 376184
rect 563568 375948 563804 376184
rect 564040 375948 564276 376184
rect 564512 375948 564748 376184
rect 564984 375948 565220 376184
rect 565456 375948 565692 376184
rect 565928 375948 566164 376184
rect 566400 375948 566636 376184
rect 566872 375948 567108 376184
rect 477192 375712 477428 375948
rect 477664 375712 477900 375948
rect 478136 375712 478372 375948
rect 478608 375712 478844 375948
rect 479080 375712 479316 375948
rect 479552 375712 479788 375948
rect 480024 375712 480260 375948
rect 480496 375712 480732 375948
rect 480968 375712 481204 375948
rect 481440 375712 481676 375948
rect 481912 375712 482148 375948
rect 482384 375712 482620 375948
rect 482856 375712 483092 375948
rect 483328 375712 483564 375948
rect 562624 375476 562860 375712
rect 563096 375476 563332 375712
rect 563568 375476 563804 375712
rect 564040 375476 564276 375712
rect 564512 375476 564748 375712
rect 564984 375476 565220 375712
rect 565456 375476 565692 375712
rect 565928 375476 566164 375712
rect 566400 375476 566636 375712
rect 566872 375476 567108 375712
rect 477192 375240 477428 375476
rect 477664 375240 477900 375476
rect 478136 375240 478372 375476
rect 478608 375240 478844 375476
rect 479080 375240 479316 375476
rect 479552 375240 479788 375476
rect 480024 375240 480260 375476
rect 480496 375240 480732 375476
rect 480968 375240 481204 375476
rect 481440 375240 481676 375476
rect 481912 375240 482148 375476
rect 482384 375240 482620 375476
rect 482856 375240 483092 375476
rect 483328 375240 483564 375476
rect 562624 375004 562860 375240
rect 563096 375004 563332 375240
rect 563568 375004 563804 375240
rect 564040 375004 564276 375240
rect 564512 375004 564748 375240
rect 564984 375004 565220 375240
rect 565456 375004 565692 375240
rect 565928 375004 566164 375240
rect 566400 375004 566636 375240
rect 566872 375004 567108 375240
rect 477192 374768 477428 375004
rect 477664 374768 477900 375004
rect 478136 374768 478372 375004
rect 478608 374768 478844 375004
rect 479080 374768 479316 375004
rect 479552 374768 479788 375004
rect 480024 374768 480260 375004
rect 480496 374768 480732 375004
rect 480968 374768 481204 375004
rect 481440 374768 481676 375004
rect 481912 374768 482148 375004
rect 482384 374768 482620 375004
rect 482856 374768 483092 375004
rect 483328 374768 483564 375004
rect 562624 374532 562860 374768
rect 563096 374532 563332 374768
rect 563568 374532 563804 374768
rect 564040 374532 564276 374768
rect 564512 374532 564748 374768
rect 564984 374532 565220 374768
rect 565456 374532 565692 374768
rect 565928 374532 566164 374768
rect 566400 374532 566636 374768
rect 566872 374532 567108 374768
rect 477192 374296 477428 374532
rect 477664 374296 477900 374532
rect 478136 374296 478372 374532
rect 478608 374296 478844 374532
rect 479080 374296 479316 374532
rect 479552 374296 479788 374532
rect 480024 374296 480260 374532
rect 480496 374296 480732 374532
rect 480968 374296 481204 374532
rect 481440 374296 481676 374532
rect 481912 374296 482148 374532
rect 482384 374296 482620 374532
rect 482856 374296 483092 374532
rect 483328 374296 483564 374532
rect 562624 374060 562860 374296
rect 563096 374060 563332 374296
rect 563568 374060 563804 374296
rect 564040 374060 564276 374296
rect 564512 374060 564748 374296
rect 564984 374060 565220 374296
rect 565456 374060 565692 374296
rect 565928 374060 566164 374296
rect 566400 374060 566636 374296
rect 566872 374060 567108 374296
rect 477192 373824 477428 374060
rect 477664 373824 477900 374060
rect 478136 373824 478372 374060
rect 478608 373824 478844 374060
rect 479080 373824 479316 374060
rect 479552 373824 479788 374060
rect 480024 373824 480260 374060
rect 480496 373824 480732 374060
rect 480968 373824 481204 374060
rect 481440 373824 481676 374060
rect 481912 373824 482148 374060
rect 482384 373824 482620 374060
rect 482856 373824 483092 374060
rect 483328 373824 483564 374060
rect 562624 373588 562860 373824
rect 563096 373588 563332 373824
rect 563568 373588 563804 373824
rect 564040 373588 564276 373824
rect 564512 373588 564748 373824
rect 564984 373588 565220 373824
rect 565456 373588 565692 373824
rect 565928 373588 566164 373824
rect 566400 373588 566636 373824
rect 566872 373588 567108 373824
rect 477192 373352 477428 373588
rect 477664 373352 477900 373588
rect 478136 373352 478372 373588
rect 478608 373352 478844 373588
rect 479080 373352 479316 373588
rect 479552 373352 479788 373588
rect 480024 373352 480260 373588
rect 480496 373352 480732 373588
rect 480968 373352 481204 373588
rect 481440 373352 481676 373588
rect 481912 373352 482148 373588
rect 482384 373352 482620 373588
rect 482856 373352 483092 373588
rect 483328 373352 483564 373588
rect 562624 373116 562860 373352
rect 563096 373116 563332 373352
rect 563568 373116 563804 373352
rect 564040 373116 564276 373352
rect 564512 373116 564748 373352
rect 564984 373116 565220 373352
rect 565456 373116 565692 373352
rect 565928 373116 566164 373352
rect 566400 373116 566636 373352
rect 566872 373116 567108 373352
rect 477192 372880 477428 373116
rect 477664 372880 477900 373116
rect 478136 372880 478372 373116
rect 478608 372880 478844 373116
rect 479080 372880 479316 373116
rect 479552 372880 479788 373116
rect 480024 372880 480260 373116
rect 480496 372880 480732 373116
rect 480968 372880 481204 373116
rect 481440 372880 481676 373116
rect 481912 372880 482148 373116
rect 482384 372880 482620 373116
rect 482856 372880 483092 373116
rect 483328 372880 483564 373116
rect 562624 372644 562860 372880
rect 563096 372644 563332 372880
rect 563568 372644 563804 372880
rect 564040 372644 564276 372880
rect 564512 372644 564748 372880
rect 564984 372644 565220 372880
rect 565456 372644 565692 372880
rect 565928 372644 566164 372880
rect 566400 372644 566636 372880
rect 566872 372644 567108 372880
rect 477192 372408 477428 372644
rect 477664 372408 477900 372644
rect 478136 372408 478372 372644
rect 478608 372408 478844 372644
rect 479080 372408 479316 372644
rect 479552 372408 479788 372644
rect 480024 372408 480260 372644
rect 480496 372408 480732 372644
rect 480968 372408 481204 372644
rect 481440 372408 481676 372644
rect 481912 372408 482148 372644
rect 482384 372408 482620 372644
rect 482856 372408 483092 372644
rect 483328 372408 483564 372644
rect 562624 372172 562860 372408
rect 563096 372172 563332 372408
rect 563568 372172 563804 372408
rect 564040 372172 564276 372408
rect 564512 372172 564748 372408
rect 564984 372172 565220 372408
rect 565456 372172 565692 372408
rect 565928 372172 566164 372408
rect 566400 372172 566636 372408
rect 566872 372172 567108 372408
rect 477192 371936 477428 372172
rect 477664 371936 477900 372172
rect 478136 371936 478372 372172
rect 478608 371936 478844 372172
rect 479080 371936 479316 372172
rect 479552 371936 479788 372172
rect 480024 371936 480260 372172
rect 480496 371936 480732 372172
rect 480968 371936 481204 372172
rect 481440 371936 481676 372172
rect 481912 371936 482148 372172
rect 482384 371936 482620 372172
rect 482856 371936 483092 372172
rect 483328 371936 483564 372172
rect 562624 371700 562860 371936
rect 563096 371700 563332 371936
rect 563568 371700 563804 371936
rect 564040 371700 564276 371936
rect 564512 371700 564748 371936
rect 564984 371700 565220 371936
rect 565456 371700 565692 371936
rect 565928 371700 566164 371936
rect 566400 371700 566636 371936
rect 566872 371700 567108 371936
rect 477192 371464 477428 371700
rect 477664 371464 477900 371700
rect 478136 371464 478372 371700
rect 478608 371464 478844 371700
rect 479080 371464 479316 371700
rect 479552 371464 479788 371700
rect 480024 371464 480260 371700
rect 480496 371464 480732 371700
rect 480968 371464 481204 371700
rect 481440 371464 481676 371700
rect 481912 371464 482148 371700
rect 482384 371464 482620 371700
rect 482856 371464 483092 371700
rect 483328 371464 483564 371700
rect 562624 371228 562860 371464
rect 563096 371228 563332 371464
rect 563568 371228 563804 371464
rect 564040 371228 564276 371464
rect 564512 371228 564748 371464
rect 564984 371228 565220 371464
rect 565456 371228 565692 371464
rect 565928 371228 566164 371464
rect 566400 371228 566636 371464
rect 566872 371228 567108 371464
<< mimcap >>
rect 511292 468700 511692 468740
rect 511292 468380 511332 468700
rect 511652 468380 511692 468700
rect 511292 468340 511692 468380
rect 511992 468700 512392 468740
rect 511992 468380 512032 468700
rect 512352 468380 512392 468700
rect 511992 468340 512392 468380
rect 512692 468700 513092 468740
rect 512692 468380 512732 468700
rect 513052 468380 513092 468700
rect 512692 468340 513092 468380
rect 513392 468700 513792 468740
rect 513392 468380 513432 468700
rect 513752 468380 513792 468700
rect 513392 468340 513792 468380
rect 514092 468700 514492 468740
rect 514092 468380 514132 468700
rect 514452 468380 514492 468700
rect 514092 468340 514492 468380
rect 514792 468700 515192 468740
rect 514792 468380 514832 468700
rect 515152 468380 515192 468700
rect 514792 468340 515192 468380
rect 515492 468700 515892 468740
rect 515492 468380 515532 468700
rect 515852 468380 515892 468700
rect 515492 468340 515892 468380
rect 516192 468700 516592 468740
rect 516192 468380 516232 468700
rect 516552 468380 516592 468700
rect 516192 468340 516592 468380
rect 516892 468700 517292 468740
rect 516892 468380 516932 468700
rect 517252 468380 517292 468700
rect 516892 468340 517292 468380
rect 517592 468700 517992 468740
rect 517592 468380 517632 468700
rect 517952 468380 517992 468700
rect 517592 468340 517992 468380
rect 511292 467981 511692 468021
rect 511292 467661 511332 467981
rect 511652 467661 511692 467981
rect 511292 467621 511692 467661
rect 511992 467981 512392 468021
rect 511992 467661 512032 467981
rect 512352 467661 512392 467981
rect 511992 467621 512392 467661
rect 512692 467981 513092 468021
rect 512692 467661 512732 467981
rect 513052 467661 513092 467981
rect 512692 467621 513092 467661
rect 513392 467981 513792 468021
rect 513392 467661 513432 467981
rect 513752 467661 513792 467981
rect 513392 467621 513792 467661
rect 514092 467981 514492 468021
rect 514092 467661 514132 467981
rect 514452 467661 514492 467981
rect 514092 467621 514492 467661
rect 514792 467981 515192 468021
rect 514792 467661 514832 467981
rect 515152 467661 515192 467981
rect 514792 467621 515192 467661
rect 515492 467981 515892 468021
rect 515492 467661 515532 467981
rect 515852 467661 515892 467981
rect 515492 467621 515892 467661
rect 516192 467981 516592 468021
rect 516192 467661 516232 467981
rect 516552 467661 516592 467981
rect 516192 467621 516592 467661
rect 516892 467981 517292 468021
rect 516892 467661 516932 467981
rect 517252 467661 517292 467981
rect 516892 467621 517292 467661
rect 517592 467981 517992 468021
rect 517592 467661 517632 467981
rect 517952 467661 517992 467981
rect 517592 467621 517992 467661
rect 511292 467262 511692 467302
rect 511292 466942 511332 467262
rect 511652 466942 511692 467262
rect 511292 466902 511692 466942
rect 511992 467262 512392 467302
rect 511992 466942 512032 467262
rect 512352 466942 512392 467262
rect 511992 466902 512392 466942
rect 512692 467262 513092 467302
rect 512692 466942 512732 467262
rect 513052 466942 513092 467262
rect 512692 466902 513092 466942
rect 513392 467262 513792 467302
rect 513392 466942 513432 467262
rect 513752 466942 513792 467262
rect 513392 466902 513792 466942
rect 514092 467262 514492 467302
rect 514092 466942 514132 467262
rect 514452 466942 514492 467262
rect 514092 466902 514492 466942
rect 514792 467262 515192 467302
rect 514792 466942 514832 467262
rect 515152 466942 515192 467262
rect 514792 466902 515192 466942
rect 515492 467262 515892 467302
rect 515492 466942 515532 467262
rect 515852 466942 515892 467262
rect 515492 466902 515892 466942
rect 516192 467262 516592 467302
rect 516192 466942 516232 467262
rect 516552 466942 516592 467262
rect 516192 466902 516592 466942
rect 516892 467262 517292 467302
rect 516892 466942 516932 467262
rect 517252 466942 517292 467262
rect 516892 466902 517292 466942
rect 517592 467262 517992 467302
rect 517592 466942 517632 467262
rect 517952 466942 517992 467262
rect 517592 466902 517992 466942
rect 511292 466543 511692 466583
rect 511292 466223 511332 466543
rect 511652 466223 511692 466543
rect 511292 466183 511692 466223
rect 511992 466543 512392 466583
rect 511992 466223 512032 466543
rect 512352 466223 512392 466543
rect 511992 466183 512392 466223
rect 512692 466543 513092 466583
rect 512692 466223 512732 466543
rect 513052 466223 513092 466543
rect 512692 466183 513092 466223
rect 513392 466543 513792 466583
rect 513392 466223 513432 466543
rect 513752 466223 513792 466543
rect 513392 466183 513792 466223
rect 514092 466543 514492 466583
rect 514092 466223 514132 466543
rect 514452 466223 514492 466543
rect 514092 466183 514492 466223
rect 514792 466543 515192 466583
rect 514792 466223 514832 466543
rect 515152 466223 515192 466543
rect 514792 466183 515192 466223
rect 515492 466543 515892 466583
rect 515492 466223 515532 466543
rect 515852 466223 515892 466543
rect 515492 466183 515892 466223
rect 516192 466543 516592 466583
rect 516192 466223 516232 466543
rect 516552 466223 516592 466543
rect 516192 466183 516592 466223
rect 516892 466543 517292 466583
rect 516892 466223 516932 466543
rect 517252 466223 517292 466543
rect 516892 466183 517292 466223
rect 517592 466543 517992 466583
rect 517592 466223 517632 466543
rect 517952 466223 517992 466543
rect 517592 466183 517992 466223
rect 511292 465824 511692 465864
rect 511292 465504 511332 465824
rect 511652 465504 511692 465824
rect 511292 465464 511692 465504
rect 511992 465824 512392 465864
rect 511992 465504 512032 465824
rect 512352 465504 512392 465824
rect 511992 465464 512392 465504
rect 512692 465824 513092 465864
rect 512692 465504 512732 465824
rect 513052 465504 513092 465824
rect 512692 465464 513092 465504
rect 513392 465824 513792 465864
rect 513392 465504 513432 465824
rect 513752 465504 513792 465824
rect 513392 465464 513792 465504
rect 514092 465824 514492 465864
rect 514092 465504 514132 465824
rect 514452 465504 514492 465824
rect 514092 465464 514492 465504
rect 514792 465824 515192 465864
rect 514792 465504 514832 465824
rect 515152 465504 515192 465824
rect 514792 465464 515192 465504
rect 515492 465824 515892 465864
rect 515492 465504 515532 465824
rect 515852 465504 515892 465824
rect 515492 465464 515892 465504
rect 516192 465824 516592 465864
rect 516192 465504 516232 465824
rect 516552 465504 516592 465824
rect 516192 465464 516592 465504
rect 516892 465824 517292 465864
rect 516892 465504 516932 465824
rect 517252 465504 517292 465824
rect 516892 465464 517292 465504
rect 517592 465824 517992 465864
rect 517592 465504 517632 465824
rect 517952 465504 517992 465824
rect 517592 465464 517992 465504
rect 511292 465105 511692 465145
rect 511292 464785 511332 465105
rect 511652 464785 511692 465105
rect 511292 464745 511692 464785
rect 511992 465105 512392 465145
rect 511992 464785 512032 465105
rect 512352 464785 512392 465105
rect 511992 464745 512392 464785
rect 512692 465105 513092 465145
rect 512692 464785 512732 465105
rect 513052 464785 513092 465105
rect 512692 464745 513092 464785
rect 513392 465105 513792 465145
rect 513392 464785 513432 465105
rect 513752 464785 513792 465105
rect 513392 464745 513792 464785
rect 514092 465105 514492 465145
rect 514092 464785 514132 465105
rect 514452 464785 514492 465105
rect 514092 464745 514492 464785
rect 514792 465105 515192 465145
rect 514792 464785 514832 465105
rect 515152 464785 515192 465105
rect 514792 464745 515192 464785
rect 515492 465105 515892 465145
rect 515492 464785 515532 465105
rect 515852 464785 515892 465105
rect 515492 464745 515892 464785
rect 516192 465105 516592 465145
rect 516192 464785 516232 465105
rect 516552 464785 516592 465105
rect 516192 464745 516592 464785
rect 516892 465105 517292 465145
rect 516892 464785 516932 465105
rect 517252 464785 517292 465105
rect 516892 464745 517292 464785
rect 517592 465105 517992 465145
rect 517592 464785 517632 465105
rect 517952 464785 517992 465105
rect 517592 464745 517992 464785
rect 511292 464386 511692 464426
rect 511292 464066 511332 464386
rect 511652 464066 511692 464386
rect 511292 464026 511692 464066
rect 511992 464386 512392 464426
rect 511992 464066 512032 464386
rect 512352 464066 512392 464386
rect 511992 464026 512392 464066
rect 512692 464386 513092 464426
rect 512692 464066 512732 464386
rect 513052 464066 513092 464386
rect 512692 464026 513092 464066
rect 513392 464386 513792 464426
rect 513392 464066 513432 464386
rect 513752 464066 513792 464386
rect 513392 464026 513792 464066
rect 514092 464386 514492 464426
rect 514092 464066 514132 464386
rect 514452 464066 514492 464386
rect 514092 464026 514492 464066
rect 514792 464386 515192 464426
rect 514792 464066 514832 464386
rect 515152 464066 515192 464386
rect 514792 464026 515192 464066
rect 515492 464386 515892 464426
rect 515492 464066 515532 464386
rect 515852 464066 515892 464386
rect 515492 464026 515892 464066
rect 516192 464386 516592 464426
rect 516192 464066 516232 464386
rect 516552 464066 516592 464386
rect 516192 464026 516592 464066
rect 516892 464386 517292 464426
rect 516892 464066 516932 464386
rect 517252 464066 517292 464386
rect 516892 464026 517292 464066
rect 517592 464386 517992 464426
rect 517592 464066 517632 464386
rect 517952 464066 517992 464386
rect 517592 464026 517992 464066
rect 511292 463667 511692 463707
rect 511292 463347 511332 463667
rect 511652 463347 511692 463667
rect 511292 463307 511692 463347
rect 511992 463667 512392 463707
rect 511992 463347 512032 463667
rect 512352 463347 512392 463667
rect 511992 463307 512392 463347
rect 512692 463667 513092 463707
rect 512692 463347 512732 463667
rect 513052 463347 513092 463667
rect 512692 463307 513092 463347
rect 513392 463667 513792 463707
rect 513392 463347 513432 463667
rect 513752 463347 513792 463667
rect 513392 463307 513792 463347
rect 514092 463667 514492 463707
rect 514092 463347 514132 463667
rect 514452 463347 514492 463667
rect 514092 463307 514492 463347
rect 514792 463667 515192 463707
rect 514792 463347 514832 463667
rect 515152 463347 515192 463667
rect 514792 463307 515192 463347
rect 515492 463667 515892 463707
rect 515492 463347 515532 463667
rect 515852 463347 515892 463667
rect 515492 463307 515892 463347
rect 516192 463667 516592 463707
rect 516192 463347 516232 463667
rect 516552 463347 516592 463667
rect 516192 463307 516592 463347
rect 516892 463667 517292 463707
rect 516892 463347 516932 463667
rect 517252 463347 517292 463667
rect 516892 463307 517292 463347
rect 517592 463667 517992 463707
rect 517592 463347 517632 463667
rect 517952 463347 517992 463667
rect 517592 463307 517992 463347
rect 511292 462948 511692 462988
rect 511292 462628 511332 462948
rect 511652 462628 511692 462948
rect 511292 462588 511692 462628
rect 511992 462948 512392 462988
rect 511992 462628 512032 462948
rect 512352 462628 512392 462948
rect 511992 462588 512392 462628
rect 512692 462948 513092 462988
rect 512692 462628 512732 462948
rect 513052 462628 513092 462948
rect 512692 462588 513092 462628
rect 513392 462948 513792 462988
rect 513392 462628 513432 462948
rect 513752 462628 513792 462948
rect 513392 462588 513792 462628
rect 514092 462948 514492 462988
rect 514092 462628 514132 462948
rect 514452 462628 514492 462948
rect 514092 462588 514492 462628
rect 514792 462948 515192 462988
rect 514792 462628 514832 462948
rect 515152 462628 515192 462948
rect 514792 462588 515192 462628
rect 515492 462948 515892 462988
rect 515492 462628 515532 462948
rect 515852 462628 515892 462948
rect 515492 462588 515892 462628
rect 516192 462948 516592 462988
rect 516192 462628 516232 462948
rect 516552 462628 516592 462948
rect 516192 462588 516592 462628
rect 516892 462948 517292 462988
rect 516892 462628 516932 462948
rect 517252 462628 517292 462948
rect 516892 462588 517292 462628
rect 517592 462948 517992 462988
rect 517592 462628 517632 462948
rect 517952 462628 517992 462948
rect 517592 462588 517992 462628
rect 511292 462229 511692 462269
rect 511292 461909 511332 462229
rect 511652 461909 511692 462229
rect 511292 461869 511692 461909
rect 511992 462229 512392 462269
rect 511992 461909 512032 462229
rect 512352 461909 512392 462229
rect 511992 461869 512392 461909
rect 512692 462229 513092 462269
rect 512692 461909 512732 462229
rect 513052 461909 513092 462229
rect 512692 461869 513092 461909
rect 513392 462229 513792 462269
rect 513392 461909 513432 462229
rect 513752 461909 513792 462229
rect 513392 461869 513792 461909
rect 514092 462229 514492 462269
rect 514092 461909 514132 462229
rect 514452 461909 514492 462229
rect 514092 461869 514492 461909
rect 514792 462229 515192 462269
rect 514792 461909 514832 462229
rect 515152 461909 515192 462229
rect 514792 461869 515192 461909
rect 515492 462229 515892 462269
rect 515492 461909 515532 462229
rect 515852 461909 515892 462229
rect 515492 461869 515892 461909
rect 516192 462229 516592 462269
rect 516192 461909 516232 462229
rect 516552 461909 516592 462229
rect 516192 461869 516592 461909
rect 516892 462229 517292 462269
rect 516892 461909 516932 462229
rect 517252 461909 517292 462229
rect 516892 461869 517292 461909
rect 517592 462229 517992 462269
rect 517592 461909 517632 462229
rect 517952 461909 517992 462229
rect 517592 461869 517992 461909
<< mimcapcontact >>
rect 511332 468380 511652 468700
rect 512032 468380 512352 468700
rect 512732 468380 513052 468700
rect 513432 468380 513752 468700
rect 514132 468380 514452 468700
rect 514832 468380 515152 468700
rect 515532 468380 515852 468700
rect 516232 468380 516552 468700
rect 516932 468380 517252 468700
rect 517632 468380 517952 468700
rect 511332 467661 511652 467981
rect 512032 467661 512352 467981
rect 512732 467661 513052 467981
rect 513432 467661 513752 467981
rect 514132 467661 514452 467981
rect 514832 467661 515152 467981
rect 515532 467661 515852 467981
rect 516232 467661 516552 467981
rect 516932 467661 517252 467981
rect 517632 467661 517952 467981
rect 511332 466942 511652 467262
rect 512032 466942 512352 467262
rect 512732 466942 513052 467262
rect 513432 466942 513752 467262
rect 514132 466942 514452 467262
rect 514832 466942 515152 467262
rect 515532 466942 515852 467262
rect 516232 466942 516552 467262
rect 516932 466942 517252 467262
rect 517632 466942 517952 467262
rect 511332 466223 511652 466543
rect 512032 466223 512352 466543
rect 512732 466223 513052 466543
rect 513432 466223 513752 466543
rect 514132 466223 514452 466543
rect 514832 466223 515152 466543
rect 515532 466223 515852 466543
rect 516232 466223 516552 466543
rect 516932 466223 517252 466543
rect 517632 466223 517952 466543
rect 511332 465504 511652 465824
rect 512032 465504 512352 465824
rect 512732 465504 513052 465824
rect 513432 465504 513752 465824
rect 514132 465504 514452 465824
rect 514832 465504 515152 465824
rect 515532 465504 515852 465824
rect 516232 465504 516552 465824
rect 516932 465504 517252 465824
rect 517632 465504 517952 465824
rect 511332 464785 511652 465105
rect 512032 464785 512352 465105
rect 512732 464785 513052 465105
rect 513432 464785 513752 465105
rect 514132 464785 514452 465105
rect 514832 464785 515152 465105
rect 515532 464785 515852 465105
rect 516232 464785 516552 465105
rect 516932 464785 517252 465105
rect 517632 464785 517952 465105
rect 511332 464066 511652 464386
rect 512032 464066 512352 464386
rect 512732 464066 513052 464386
rect 513432 464066 513752 464386
rect 514132 464066 514452 464386
rect 514832 464066 515152 464386
rect 515532 464066 515852 464386
rect 516232 464066 516552 464386
rect 516932 464066 517252 464386
rect 517632 464066 517952 464386
rect 511332 463347 511652 463667
rect 512032 463347 512352 463667
rect 512732 463347 513052 463667
rect 513432 463347 513752 463667
rect 514132 463347 514452 463667
rect 514832 463347 515152 463667
rect 515532 463347 515852 463667
rect 516232 463347 516552 463667
rect 516932 463347 517252 463667
rect 517632 463347 517952 463667
rect 511332 462628 511652 462948
rect 512032 462628 512352 462948
rect 512732 462628 513052 462948
rect 513432 462628 513752 462948
rect 514132 462628 514452 462948
rect 514832 462628 515152 462948
rect 515532 462628 515852 462948
rect 516232 462628 516552 462948
rect 516932 462628 517252 462948
rect 517632 462628 517952 462948
rect 511332 461909 511652 462229
rect 512032 461909 512352 462229
rect 512732 461909 513052 462229
rect 513432 461909 513752 462229
rect 514132 461909 514452 462229
rect 514832 461909 515152 462229
rect 515532 461909 515852 462229
rect 516232 461909 516552 462229
rect 516932 461909 517252 462229
rect 517632 461909 517952 462229
<< metal4 >>
rect 115334 697380 577480 697420
rect 115334 697360 577492 697380
rect 115334 697200 510654 697360
rect 115334 692600 171000 697200
rect 173000 692600 173400 697200
rect 175400 692600 222706 697200
rect 224706 692600 225106 697200
rect 227106 692600 324412 697200
rect 326412 692600 326812 697200
rect 328812 692600 510654 697200
rect 115334 692560 510654 692600
rect 515334 692560 520654 697360
rect 525334 697144 577492 697360
rect 525334 696908 572772 697144
rect 573008 696908 573244 697144
rect 573480 696908 573716 697144
rect 573952 696908 574188 697144
rect 574424 696908 574660 697144
rect 574896 696908 575132 697144
rect 575368 696908 575604 697144
rect 575840 696908 576076 697144
rect 576312 696908 576548 697144
rect 576784 696908 577020 697144
rect 577256 696908 577492 697144
rect 525334 696672 577492 696908
rect 525334 696436 572772 696672
rect 573008 696436 573244 696672
rect 573480 696436 573716 696672
rect 573952 696436 574188 696672
rect 574424 696436 574660 696672
rect 574896 696436 575132 696672
rect 575368 696436 575604 696672
rect 575840 696436 576076 696672
rect 576312 696436 576548 696672
rect 576784 696436 577020 696672
rect 577256 696436 577492 696672
rect 525334 696200 577492 696436
rect 525334 695964 572772 696200
rect 573008 695964 573244 696200
rect 573480 695964 573716 696200
rect 573952 695964 574188 696200
rect 574424 695964 574660 696200
rect 574896 695964 575132 696200
rect 575368 695964 575604 696200
rect 575840 695964 576076 696200
rect 576312 695964 576548 696200
rect 576784 695964 577020 696200
rect 577256 695964 577492 696200
rect 525334 695728 577492 695964
rect 525334 695492 572772 695728
rect 573008 695492 573244 695728
rect 573480 695492 573716 695728
rect 573952 695492 574188 695728
rect 574424 695492 574660 695728
rect 574896 695492 575132 695728
rect 575368 695492 575604 695728
rect 575840 695492 576076 695728
rect 576312 695492 576548 695728
rect 576784 695492 577020 695728
rect 577256 695492 577492 695728
rect 525334 695256 577492 695492
rect 525334 695020 572772 695256
rect 573008 695020 573244 695256
rect 573480 695020 573716 695256
rect 573952 695020 574188 695256
rect 574424 695020 574660 695256
rect 574896 695020 575132 695256
rect 575368 695020 575604 695256
rect 575840 695020 576076 695256
rect 576312 695020 576548 695256
rect 576784 695020 577020 695256
rect 577256 695020 577492 695256
rect 525334 694784 577492 695020
rect 525334 694548 572772 694784
rect 573008 694548 573244 694784
rect 573480 694548 573716 694784
rect 573952 694548 574188 694784
rect 574424 694548 574660 694784
rect 574896 694548 575132 694784
rect 575368 694548 575604 694784
rect 575840 694548 576076 694784
rect 576312 694548 576548 694784
rect 576784 694548 577020 694784
rect 577256 694548 577492 694784
rect 525334 694312 577492 694548
rect 525334 694076 572772 694312
rect 573008 694076 573244 694312
rect 573480 694076 573716 694312
rect 573952 694076 574188 694312
rect 574424 694076 574660 694312
rect 574896 694076 575132 694312
rect 575368 694076 575604 694312
rect 575840 694076 576076 694312
rect 576312 694076 576548 694312
rect 576784 694076 577020 694312
rect 577256 694076 577492 694312
rect 525334 693840 577492 694076
rect 525334 693604 572772 693840
rect 573008 693604 573244 693840
rect 573480 693604 573716 693840
rect 573952 693604 574188 693840
rect 574424 693604 574660 693840
rect 574896 693604 575132 693840
rect 575368 693604 575604 693840
rect 575840 693604 576076 693840
rect 576312 693604 576548 693840
rect 576784 693604 577020 693840
rect 577256 693604 577492 693840
rect 525334 693368 577492 693604
rect 525334 693132 572772 693368
rect 573008 693132 573244 693368
rect 573480 693132 573716 693368
rect 573952 693132 574188 693368
rect 574424 693132 574660 693368
rect 574896 693132 575132 693368
rect 575368 693132 575604 693368
rect 575840 693132 576076 693368
rect 576312 693132 576548 693368
rect 576784 693132 577020 693368
rect 577256 693132 577492 693368
rect 525334 692896 577492 693132
rect 525334 692660 572772 692896
rect 573008 692660 573244 692896
rect 573480 692660 573716 692896
rect 573952 692660 574188 692896
rect 574424 692660 574660 692896
rect 574896 692660 575132 692896
rect 575368 692660 575604 692896
rect 575840 692660 576076 692896
rect 576312 692660 576548 692896
rect 576784 692660 577020 692896
rect 577256 692660 577492 692896
rect 525334 692560 577480 692660
rect 115334 692500 577480 692560
rect 562456 644584 567424 644608
rect 562456 639784 562480 644584
rect 567400 639784 567424 644584
rect 562456 639760 567424 639784
rect 562456 634584 567424 634608
rect 562456 629784 562480 634584
rect 567400 629784 567424 634584
rect 562456 629760 567424 629784
rect 572600 623400 577400 623588
rect 477192 522892 483800 523098
rect 477060 522862 483800 522892
rect 477060 522626 477192 522862
rect 477428 522626 477664 522862
rect 477900 522626 478136 522862
rect 478372 522626 478608 522862
rect 478844 522626 479080 522862
rect 479316 522626 479552 522862
rect 479788 522626 480024 522862
rect 480260 522626 480496 522862
rect 480732 522626 480968 522862
rect 481204 522626 481440 522862
rect 481676 522626 481912 522862
rect 482148 522626 482384 522862
rect 482620 522626 482856 522862
rect 483092 522626 483328 522862
rect 483564 522626 483800 522862
rect 477060 522390 483800 522626
rect 477060 522154 477192 522390
rect 477428 522154 477664 522390
rect 477900 522154 478136 522390
rect 478372 522154 478608 522390
rect 478844 522154 479080 522390
rect 479316 522154 479552 522390
rect 479788 522154 480024 522390
rect 480260 522154 480496 522390
rect 480732 522154 480968 522390
rect 481204 522154 481440 522390
rect 481676 522154 481912 522390
rect 482148 522154 482384 522390
rect 482620 522154 482856 522390
rect 483092 522154 483328 522390
rect 483564 522154 483800 522390
rect 477060 521918 483800 522154
rect 477060 521682 477192 521918
rect 477428 521682 477664 521918
rect 477900 521682 478136 521918
rect 478372 521682 478608 521918
rect 478844 521682 479080 521918
rect 479316 521682 479552 521918
rect 479788 521682 480024 521918
rect 480260 521682 480496 521918
rect 480732 521682 480968 521918
rect 481204 521682 481440 521918
rect 481676 521682 481912 521918
rect 482148 521682 482384 521918
rect 482620 521682 482856 521918
rect 483092 521682 483328 521918
rect 483564 521682 483800 521918
rect 477060 521446 483800 521682
rect 477060 521210 477192 521446
rect 477428 521210 477664 521446
rect 477900 521210 478136 521446
rect 478372 521210 478608 521446
rect 478844 521210 479080 521446
rect 479316 521210 479552 521446
rect 479788 521210 480024 521446
rect 480260 521210 480496 521446
rect 480732 521210 480968 521446
rect 481204 521210 481440 521446
rect 481676 521210 481912 521446
rect 482148 521210 482384 521446
rect 482620 521210 482856 521446
rect 483092 521210 483328 521446
rect 483564 521210 483800 521446
rect 477060 520974 483800 521210
rect 477060 520738 477192 520974
rect 477428 520738 477664 520974
rect 477900 520738 478136 520974
rect 478372 520738 478608 520974
rect 478844 520738 479080 520974
rect 479316 520738 479552 520974
rect 479788 520738 480024 520974
rect 480260 520738 480496 520974
rect 480732 520738 480968 520974
rect 481204 520738 481440 520974
rect 481676 520738 481912 520974
rect 482148 520738 482384 520974
rect 482620 520738 482856 520974
rect 483092 520738 483328 520974
rect 483564 520738 483800 520974
rect 477060 520502 483800 520738
rect 477060 520266 477192 520502
rect 477428 520266 477664 520502
rect 477900 520266 478136 520502
rect 478372 520266 478608 520502
rect 478844 520266 479080 520502
rect 479316 520266 479552 520502
rect 479788 520266 480024 520502
rect 480260 520266 480496 520502
rect 480732 520266 480968 520502
rect 481204 520266 481440 520502
rect 481676 520266 481912 520502
rect 482148 520266 482384 520502
rect 482620 520266 482856 520502
rect 483092 520266 483328 520502
rect 483564 520266 483800 520502
rect 477060 520030 483800 520266
rect 477060 519794 477192 520030
rect 477428 519794 477664 520030
rect 477900 519794 478136 520030
rect 478372 519794 478608 520030
rect 478844 519794 479080 520030
rect 479316 519794 479552 520030
rect 479788 519794 480024 520030
rect 480260 519794 480496 520030
rect 480732 519794 480968 520030
rect 481204 519794 481440 520030
rect 481676 519794 481912 520030
rect 482148 519794 482384 520030
rect 482620 519794 482856 520030
rect 483092 519794 483328 520030
rect 483564 519794 483800 520030
rect 477060 519558 483800 519794
rect 477060 519322 477192 519558
rect 477428 519322 477664 519558
rect 477900 519322 478136 519558
rect 478372 519322 478608 519558
rect 478844 519322 479080 519558
rect 479316 519322 479552 519558
rect 479788 519322 480024 519558
rect 480260 519322 480496 519558
rect 480732 519322 480968 519558
rect 481204 519322 481440 519558
rect 481676 519322 481912 519558
rect 482148 519322 482384 519558
rect 482620 519322 482856 519558
rect 483092 519322 483328 519558
rect 483564 519322 483800 519558
rect 477060 519086 483800 519322
rect 477060 518850 477192 519086
rect 477428 518850 477664 519086
rect 477900 518850 478136 519086
rect 478372 518850 478608 519086
rect 478844 518850 479080 519086
rect 479316 518850 479552 519086
rect 479788 518850 480024 519086
rect 480260 518850 480496 519086
rect 480732 518850 480968 519086
rect 481204 518850 481440 519086
rect 481676 518850 481912 519086
rect 482148 518850 482384 519086
rect 482620 518850 482856 519086
rect 483092 518850 483328 519086
rect 483564 518850 483800 519086
rect 477060 518614 483800 518850
rect 477060 518378 477192 518614
rect 477428 518378 477664 518614
rect 477900 518378 478136 518614
rect 478372 518378 478608 518614
rect 478844 518378 479080 518614
rect 479316 518378 479552 518614
rect 479788 518378 480024 518614
rect 480260 518378 480496 518614
rect 480732 518378 480968 518614
rect 481204 518378 481440 518614
rect 481676 518378 481912 518614
rect 482148 518378 482384 518614
rect 482620 518378 482856 518614
rect 483092 518378 483328 518614
rect 483564 518378 483800 518614
rect 477060 518142 483800 518378
rect 477060 517906 477192 518142
rect 477428 517906 477664 518142
rect 477900 517906 478136 518142
rect 478372 517906 478608 518142
rect 478844 517906 479080 518142
rect 479316 517906 479552 518142
rect 479788 517906 480024 518142
rect 480260 517906 480496 518142
rect 480732 517906 480968 518142
rect 481204 517906 481440 518142
rect 481676 517906 481912 518142
rect 482148 517906 482384 518142
rect 482620 517906 482856 518142
rect 483092 517906 483328 518142
rect 483564 517906 483800 518142
rect 477060 517670 483800 517906
rect 477060 517434 477192 517670
rect 477428 517434 477664 517670
rect 477900 517434 478136 517670
rect 478372 517434 478608 517670
rect 478844 517434 479080 517670
rect 479316 517434 479552 517670
rect 479788 517434 480024 517670
rect 480260 517434 480496 517670
rect 480732 517434 480968 517670
rect 481204 517434 481440 517670
rect 481676 517434 481912 517670
rect 482148 517434 482384 517670
rect 482620 517434 482856 517670
rect 483092 517434 483328 517670
rect 483564 517434 483800 517670
rect 477060 517198 483800 517434
rect 477060 516962 477192 517198
rect 477428 516962 477664 517198
rect 477900 516962 478136 517198
rect 478372 516962 478608 517198
rect 478844 516962 479080 517198
rect 479316 516962 479552 517198
rect 479788 516962 480024 517198
rect 480260 516962 480496 517198
rect 480732 516962 480968 517198
rect 481204 516962 481440 517198
rect 481676 516962 481912 517198
rect 482148 516962 482384 517198
rect 482620 516962 482856 517198
rect 483092 516962 483328 517198
rect 483564 516962 483800 517198
rect 477060 516726 483800 516962
rect 477060 516490 477192 516726
rect 477428 516490 477664 516726
rect 477900 516490 478136 516726
rect 478372 516490 478608 516726
rect 478844 516490 479080 516726
rect 479316 516490 479552 516726
rect 479788 516490 480024 516726
rect 480260 516490 480496 516726
rect 480732 516490 480968 516726
rect 481204 516490 481440 516726
rect 481676 516490 481912 516726
rect 482148 516490 482384 516726
rect 482620 516490 482856 516726
rect 483092 516490 483328 516726
rect 483564 516490 483800 516726
rect 562388 522740 567816 523212
rect 477060 455676 483726 516490
rect 562388 516368 562624 522740
rect 562860 516368 563096 522740
rect 563332 516368 563568 522740
rect 563804 516368 564040 522740
rect 564276 516368 564512 522740
rect 564748 516368 564984 522740
rect 565220 516368 565456 522740
rect 565692 516368 565928 522740
rect 566164 516368 566400 522740
rect 566636 516368 566872 522740
rect 567108 516368 567816 522740
rect 562388 516132 567816 516368
rect 562380 495782 567480 495822
rect 562380 495742 562624 495782
rect 562860 495742 563096 495782
rect 563332 495742 563568 495782
rect 563804 495742 564040 495782
rect 564276 495742 564512 495782
rect 564748 495742 564984 495782
rect 565220 495742 565456 495782
rect 565692 495742 565928 495782
rect 566164 495742 566400 495782
rect 566636 495742 566872 495782
rect 567108 495742 567480 495782
rect 562380 495662 562480 495742
rect 562560 495662 562624 495742
rect 562880 495662 562960 495742
rect 563040 495662 563096 495742
rect 563360 495662 563440 495742
rect 563520 495662 563568 495742
rect 563840 495662 563920 495742
rect 564000 495662 564040 495742
rect 564320 495662 564400 495742
rect 564480 495662 564512 495742
rect 564800 495662 564880 495742
rect 564960 495662 564984 495742
rect 565280 495662 565360 495742
rect 565440 495662 565456 495742
rect 565760 495662 565840 495742
rect 565920 495662 565928 495742
rect 566240 495662 566320 495742
rect 566636 495662 566640 495742
rect 566720 495662 566800 495742
rect 567108 495662 567120 495742
rect 567200 495662 567280 495742
rect 567360 495662 567480 495742
rect 562380 495582 562624 495662
rect 562860 495582 563096 495662
rect 563332 495582 563568 495662
rect 563804 495582 564040 495662
rect 564276 495582 564512 495662
rect 564748 495582 564984 495662
rect 565220 495582 565456 495662
rect 565692 495582 565928 495662
rect 566164 495582 566400 495662
rect 566636 495582 566872 495662
rect 567108 495582 567480 495662
rect 562380 495502 562480 495582
rect 562560 495546 562624 495582
rect 562560 495502 562640 495546
rect 562720 495502 562800 495546
rect 562880 495502 562960 495582
rect 563040 495546 563096 495582
rect 563040 495502 563120 495546
rect 563200 495502 563280 495546
rect 563360 495502 563440 495582
rect 563520 495546 563568 495582
rect 563520 495502 563600 495546
rect 563680 495502 563760 495546
rect 563840 495502 563920 495582
rect 564000 495546 564040 495582
rect 564000 495502 564080 495546
rect 564160 495502 564240 495546
rect 564320 495502 564400 495582
rect 564480 495546 564512 495582
rect 564480 495502 564560 495546
rect 564640 495502 564720 495546
rect 564800 495502 564880 495582
rect 564960 495546 564984 495582
rect 564960 495502 565040 495546
rect 565120 495502 565200 495546
rect 565280 495502 565360 495582
rect 565440 495546 565456 495582
rect 565440 495502 565520 495546
rect 565600 495502 565680 495546
rect 565760 495502 565840 495582
rect 565920 495546 565928 495582
rect 565920 495502 566000 495546
rect 566080 495502 566160 495546
rect 566240 495502 566320 495582
rect 566636 495546 566640 495582
rect 566400 495502 566480 495546
rect 566560 495502 566640 495546
rect 566720 495502 566800 495582
rect 567108 495546 567120 495582
rect 566880 495502 566960 495546
rect 567040 495502 567120 495546
rect 567200 495502 567280 495582
rect 567360 495502 567480 495582
rect 562380 495462 567480 495502
rect 572540 495782 577640 495822
rect 572540 495742 572784 495782
rect 573020 495742 573256 495782
rect 573492 495742 573728 495782
rect 573964 495742 574200 495782
rect 574436 495742 574672 495782
rect 574908 495742 575144 495782
rect 575380 495742 575616 495782
rect 575852 495742 576088 495782
rect 576324 495742 576560 495782
rect 576796 495742 577032 495782
rect 577268 495742 577640 495782
rect 572540 495662 572640 495742
rect 572720 495662 572784 495742
rect 573040 495662 573120 495742
rect 573200 495662 573256 495742
rect 573520 495662 573600 495742
rect 573680 495662 573728 495742
rect 574000 495662 574080 495742
rect 574160 495662 574200 495742
rect 574480 495662 574560 495742
rect 574640 495662 574672 495742
rect 574960 495662 575040 495742
rect 575120 495662 575144 495742
rect 575440 495662 575520 495742
rect 575600 495662 575616 495742
rect 575920 495662 576000 495742
rect 576080 495662 576088 495742
rect 576400 495662 576480 495742
rect 576796 495662 576800 495742
rect 576880 495662 576960 495742
rect 577268 495662 577280 495742
rect 577360 495662 577440 495742
rect 577520 495662 577640 495742
rect 572540 495582 572784 495662
rect 573020 495582 573256 495662
rect 573492 495582 573728 495662
rect 573964 495582 574200 495662
rect 574436 495582 574672 495662
rect 574908 495582 575144 495662
rect 575380 495582 575616 495662
rect 575852 495582 576088 495662
rect 576324 495582 576560 495662
rect 576796 495582 577032 495662
rect 577268 495582 577640 495662
rect 572540 495502 572640 495582
rect 572720 495546 572784 495582
rect 572720 495502 572800 495546
rect 572880 495502 572960 495546
rect 573040 495502 573120 495582
rect 573200 495546 573256 495582
rect 573200 495502 573280 495546
rect 573360 495502 573440 495546
rect 573520 495502 573600 495582
rect 573680 495546 573728 495582
rect 573680 495502 573760 495546
rect 573840 495502 573920 495546
rect 574000 495502 574080 495582
rect 574160 495546 574200 495582
rect 574160 495502 574240 495546
rect 574320 495502 574400 495546
rect 574480 495502 574560 495582
rect 574640 495546 574672 495582
rect 574640 495502 574720 495546
rect 574800 495502 574880 495546
rect 574960 495502 575040 495582
rect 575120 495546 575144 495582
rect 575120 495502 575200 495546
rect 575280 495502 575360 495546
rect 575440 495502 575520 495582
rect 575600 495546 575616 495582
rect 575600 495502 575680 495546
rect 575760 495502 575840 495546
rect 575920 495502 576000 495582
rect 576080 495546 576088 495582
rect 576080 495502 576160 495546
rect 576240 495502 576320 495546
rect 576400 495502 576480 495582
rect 576796 495546 576800 495582
rect 576560 495502 576640 495546
rect 576720 495502 576800 495546
rect 576880 495502 576960 495582
rect 577268 495546 577280 495582
rect 577040 495502 577120 495546
rect 577200 495502 577280 495546
rect 577360 495502 577440 495582
rect 577520 495502 577640 495582
rect 572540 495462 577640 495502
rect 511584 494528 512160 494700
rect 511584 494464 511616 494528
rect 511680 494464 511744 494528
rect 511808 494464 511872 494528
rect 511936 494464 512000 494528
rect 512064 494464 512160 494528
rect 511584 494400 512160 494464
rect 511584 494336 511616 494400
rect 511680 494336 511744 494400
rect 511808 494336 511872 494400
rect 511936 494336 512000 494400
rect 512064 494336 512160 494400
rect 511584 494272 512160 494336
rect 511584 494208 511616 494272
rect 511680 494208 511744 494272
rect 511808 494208 511872 494272
rect 511936 494208 512000 494272
rect 512064 494208 512160 494272
rect 511584 494144 512160 494208
rect 511584 494080 511616 494144
rect 511680 494080 511744 494144
rect 511808 494080 511872 494144
rect 511936 494080 512000 494144
rect 512064 494080 512160 494144
rect 511584 494016 512160 494080
rect 511584 493952 511616 494016
rect 511680 493952 511744 494016
rect 511808 493952 511872 494016
rect 511936 493952 512000 494016
rect 512064 493952 512160 494016
rect 511584 493888 512160 493952
rect 511584 493824 511616 493888
rect 511680 493824 511744 493888
rect 511808 493824 511872 493888
rect 511936 493824 512000 493888
rect 512064 493824 512160 493888
rect 490440 483236 497096 487356
rect 490440 478452 490940 483236
rect 496684 478452 497096 483236
rect 490440 474236 497096 478452
rect 503860 483236 510540 484136
rect 503860 478452 503960 483236
rect 509704 478452 510540 483236
rect 503860 475306 510540 478452
rect 503860 475206 503920 475306
rect 504020 475206 504144 475306
rect 504244 475206 504368 475306
rect 504468 475206 504592 475306
rect 504692 475206 504816 475306
rect 504916 475206 505040 475306
rect 505140 475206 505264 475306
rect 505364 475206 505488 475306
rect 505588 475206 505712 475306
rect 505812 475206 505936 475306
rect 506036 475206 506160 475306
rect 506260 475206 506384 475306
rect 506484 475206 506608 475306
rect 506708 475206 506832 475306
rect 506932 475206 507056 475306
rect 507156 475206 507280 475306
rect 507380 475206 507504 475306
rect 507604 475206 507728 475306
rect 507828 475206 507952 475306
rect 508052 475206 508176 475306
rect 508276 475206 508400 475306
rect 508500 475206 508624 475306
rect 508724 475206 508848 475306
rect 508948 475206 509072 475306
rect 509172 475206 509296 475306
rect 509396 475206 509520 475306
rect 509620 475206 509744 475306
rect 509844 475206 509968 475306
rect 510068 475206 510192 475306
rect 510292 475206 510416 475306
rect 510516 475206 510540 475306
rect 503860 475082 510540 475206
rect 503860 474982 503920 475082
rect 504020 474982 504144 475082
rect 504244 474982 504368 475082
rect 504468 474982 504592 475082
rect 504692 474982 504816 475082
rect 504916 474982 505040 475082
rect 505140 474982 505264 475082
rect 505364 474982 505488 475082
rect 505588 474982 505712 475082
rect 505812 474982 505936 475082
rect 506036 474982 506160 475082
rect 506260 474982 506384 475082
rect 506484 474982 506608 475082
rect 506708 474982 506832 475082
rect 506932 474982 507056 475082
rect 507156 474982 507280 475082
rect 507380 474982 507504 475082
rect 507604 474982 507728 475082
rect 507828 474982 507952 475082
rect 508052 474982 508176 475082
rect 508276 474982 508400 475082
rect 508500 474982 508624 475082
rect 508724 474982 508848 475082
rect 508948 474982 509072 475082
rect 509172 474982 509296 475082
rect 509396 474982 509520 475082
rect 509620 474982 509744 475082
rect 509844 474982 509968 475082
rect 510068 474982 510192 475082
rect 510292 474982 510416 475082
rect 510516 474982 510540 475082
rect 503860 474858 510540 474982
rect 503860 474758 503920 474858
rect 504020 474758 504144 474858
rect 504244 474758 504368 474858
rect 504468 474758 504592 474858
rect 504692 474758 504816 474858
rect 504916 474758 505040 474858
rect 505140 474758 505264 474858
rect 505364 474758 505488 474858
rect 505588 474758 505712 474858
rect 505812 474758 505936 474858
rect 506036 474758 506160 474858
rect 506260 474758 506384 474858
rect 506484 474758 506608 474858
rect 506708 474758 506832 474858
rect 506932 474758 507056 474858
rect 507156 474758 507280 474858
rect 507380 474758 507504 474858
rect 507604 474758 507728 474858
rect 507828 474758 507952 474858
rect 508052 474758 508176 474858
rect 508276 474758 508400 474858
rect 508500 474758 508624 474858
rect 508724 474758 508848 474858
rect 508948 474758 509072 474858
rect 509172 474758 509296 474858
rect 509396 474758 509520 474858
rect 509620 474758 509744 474858
rect 509844 474758 509968 474858
rect 510068 474758 510192 474858
rect 510292 474758 510416 474858
rect 510516 474758 510540 474858
rect 503860 474634 510540 474758
rect 503860 474534 503920 474634
rect 504020 474534 504144 474634
rect 504244 474534 504368 474634
rect 504468 474534 504592 474634
rect 504692 474534 504816 474634
rect 504916 474534 505040 474634
rect 505140 474534 505264 474634
rect 505364 474534 505488 474634
rect 505588 474534 505712 474634
rect 505812 474534 505936 474634
rect 506036 474534 506160 474634
rect 506260 474534 506384 474634
rect 506484 474534 506608 474634
rect 506708 474534 506832 474634
rect 506932 474534 507056 474634
rect 507156 474534 507280 474634
rect 507380 474534 507504 474634
rect 507604 474534 507728 474634
rect 507828 474534 507952 474634
rect 508052 474534 508176 474634
rect 508276 474534 508400 474634
rect 508500 474534 508624 474634
rect 508724 474534 508848 474634
rect 508948 474534 509072 474634
rect 509172 474534 509296 474634
rect 509396 474534 509520 474634
rect 509620 474534 509744 474634
rect 509844 474534 509968 474634
rect 510068 474534 510192 474634
rect 510292 474534 510416 474634
rect 510516 474534 510540 474634
rect 503860 474410 510540 474534
rect 490440 469452 491256 474236
rect 497000 469452 497096 474236
rect 490440 468236 497096 469452
rect 490440 463452 491256 468236
rect 497000 463452 497096 468236
rect 500364 474280 501404 474336
rect 500364 474180 500398 474280
rect 500498 474180 500622 474280
rect 500722 474180 500846 474280
rect 500946 474180 501070 474280
rect 501170 474180 501294 474280
rect 501394 474180 501404 474280
rect 503860 474310 503920 474410
rect 504020 474310 504144 474410
rect 504244 474310 504368 474410
rect 504468 474310 504592 474410
rect 504692 474310 504816 474410
rect 504916 474310 505040 474410
rect 505140 474310 505264 474410
rect 505364 474310 505488 474410
rect 505588 474310 505712 474410
rect 505812 474310 505936 474410
rect 506036 474310 506160 474410
rect 506260 474310 506384 474410
rect 506484 474310 506608 474410
rect 506708 474310 506832 474410
rect 506932 474310 507056 474410
rect 507156 474310 507280 474410
rect 507380 474310 507504 474410
rect 507604 474310 507728 474410
rect 507828 474310 507952 474410
rect 508052 474310 508176 474410
rect 508276 474310 508400 474410
rect 508500 474310 508624 474410
rect 508724 474310 508848 474410
rect 508948 474310 509072 474410
rect 509172 474310 509296 474410
rect 509396 474310 509520 474410
rect 509620 474310 509744 474410
rect 509844 474310 509968 474410
rect 510068 474310 510192 474410
rect 510292 474310 510416 474410
rect 510516 474310 510540 474410
rect 503860 474276 510540 474310
rect 511584 475300 512160 493824
rect 511584 475236 511648 475300
rect 511712 475236 511776 475300
rect 511840 475236 511904 475300
rect 511968 475236 512032 475300
rect 512096 475236 512160 475300
rect 511584 475172 512160 475236
rect 511584 475108 511648 475172
rect 511712 475108 511776 475172
rect 511840 475108 511904 475172
rect 511968 475108 512032 475172
rect 512096 475108 512160 475172
rect 511584 475044 512160 475108
rect 511584 474980 511648 475044
rect 511712 474980 511776 475044
rect 511840 474980 511904 475044
rect 511968 474980 512032 475044
rect 512096 474980 512160 475044
rect 511584 474916 512160 474980
rect 511584 474852 511648 474916
rect 511712 474852 511776 474916
rect 511840 474852 511904 474916
rect 511968 474852 512032 474916
rect 512096 474852 512160 474916
rect 511584 474788 512160 474852
rect 511584 474724 511648 474788
rect 511712 474724 511776 474788
rect 511840 474724 511904 474788
rect 511968 474724 512032 474788
rect 512096 474724 512160 474788
rect 511584 474660 512160 474724
rect 511584 474596 511648 474660
rect 511712 474596 511776 474660
rect 511840 474596 511904 474660
rect 511968 474596 512032 474660
rect 512096 474596 512160 474660
rect 511584 474532 512160 474596
rect 511584 474468 511648 474532
rect 511712 474468 511776 474532
rect 511840 474468 511904 474532
rect 511968 474468 512032 474532
rect 512096 474468 512160 474532
rect 511584 474404 512160 474468
rect 511584 474340 511648 474404
rect 511712 474340 511776 474404
rect 511840 474340 511904 474404
rect 511968 474340 512032 474404
rect 512096 474340 512160 474404
rect 511584 474276 512160 474340
rect 517260 483236 523940 484136
rect 517260 478452 517360 483236
rect 523104 478452 523940 483236
rect 517260 475306 523940 478452
rect 517260 475206 517320 475306
rect 517420 475206 517544 475306
rect 517644 475206 517768 475306
rect 517868 475206 517992 475306
rect 518092 475206 518216 475306
rect 518316 475206 518440 475306
rect 518540 475206 518664 475306
rect 518764 475206 518888 475306
rect 518988 475206 519112 475306
rect 519212 475206 519336 475306
rect 519436 475206 519560 475306
rect 519660 475206 519784 475306
rect 519884 475206 520008 475306
rect 520108 475206 520232 475306
rect 520332 475206 520456 475306
rect 520556 475206 520680 475306
rect 520780 475206 520904 475306
rect 521004 475206 521128 475306
rect 521228 475206 521352 475306
rect 521452 475206 521576 475306
rect 521676 475206 521800 475306
rect 521900 475206 522024 475306
rect 522124 475206 522248 475306
rect 522348 475206 522472 475306
rect 522572 475206 522696 475306
rect 522796 475206 522920 475306
rect 523020 475206 523144 475306
rect 523244 475206 523368 475306
rect 523468 475206 523592 475306
rect 523692 475206 523816 475306
rect 523916 475206 523940 475306
rect 517260 475082 523940 475206
rect 517260 474982 517320 475082
rect 517420 474982 517544 475082
rect 517644 474982 517768 475082
rect 517868 474982 517992 475082
rect 518092 474982 518216 475082
rect 518316 474982 518440 475082
rect 518540 474982 518664 475082
rect 518764 474982 518888 475082
rect 518988 474982 519112 475082
rect 519212 474982 519336 475082
rect 519436 474982 519560 475082
rect 519660 474982 519784 475082
rect 519884 474982 520008 475082
rect 520108 474982 520232 475082
rect 520332 474982 520456 475082
rect 520556 474982 520680 475082
rect 520780 474982 520904 475082
rect 521004 474982 521128 475082
rect 521228 474982 521352 475082
rect 521452 474982 521576 475082
rect 521676 474982 521800 475082
rect 521900 474982 522024 475082
rect 522124 474982 522248 475082
rect 522348 474982 522472 475082
rect 522572 474982 522696 475082
rect 522796 474982 522920 475082
rect 523020 474982 523144 475082
rect 523244 474982 523368 475082
rect 523468 474982 523592 475082
rect 523692 474982 523816 475082
rect 523916 474982 523940 475082
rect 517260 474858 523940 474982
rect 517260 474758 517320 474858
rect 517420 474758 517544 474858
rect 517644 474758 517768 474858
rect 517868 474758 517992 474858
rect 518092 474758 518216 474858
rect 518316 474758 518440 474858
rect 518540 474758 518664 474858
rect 518764 474758 518888 474858
rect 518988 474758 519112 474858
rect 519212 474758 519336 474858
rect 519436 474758 519560 474858
rect 519660 474758 519784 474858
rect 519884 474758 520008 474858
rect 520108 474758 520232 474858
rect 520332 474758 520456 474858
rect 520556 474758 520680 474858
rect 520780 474758 520904 474858
rect 521004 474758 521128 474858
rect 521228 474758 521352 474858
rect 521452 474758 521576 474858
rect 521676 474758 521800 474858
rect 521900 474758 522024 474858
rect 522124 474758 522248 474858
rect 522348 474758 522472 474858
rect 522572 474758 522696 474858
rect 522796 474758 522920 474858
rect 523020 474758 523144 474858
rect 523244 474758 523368 474858
rect 523468 474758 523592 474858
rect 523692 474758 523816 474858
rect 523916 474758 523940 474858
rect 517260 474634 523940 474758
rect 517260 474534 517320 474634
rect 517420 474534 517544 474634
rect 517644 474534 517768 474634
rect 517868 474534 517992 474634
rect 518092 474534 518216 474634
rect 518316 474534 518440 474634
rect 518540 474534 518664 474634
rect 518764 474534 518888 474634
rect 518988 474534 519112 474634
rect 519212 474534 519336 474634
rect 519436 474534 519560 474634
rect 519660 474534 519784 474634
rect 519884 474534 520008 474634
rect 520108 474534 520232 474634
rect 520332 474534 520456 474634
rect 520556 474534 520680 474634
rect 520780 474534 520904 474634
rect 521004 474534 521128 474634
rect 521228 474534 521352 474634
rect 521452 474534 521576 474634
rect 521676 474534 521800 474634
rect 521900 474534 522024 474634
rect 522124 474534 522248 474634
rect 522348 474534 522472 474634
rect 522572 474534 522696 474634
rect 522796 474534 522920 474634
rect 523020 474534 523144 474634
rect 523244 474534 523368 474634
rect 523468 474534 523592 474634
rect 523692 474534 523816 474634
rect 523916 474534 523940 474634
rect 517260 474410 523940 474534
rect 517260 474310 517320 474410
rect 517420 474310 517544 474410
rect 517644 474310 517768 474410
rect 517868 474310 517992 474410
rect 518092 474310 518216 474410
rect 518316 474310 518440 474410
rect 518540 474310 518664 474410
rect 518764 474310 518888 474410
rect 518988 474310 519112 474410
rect 519212 474310 519336 474410
rect 519436 474310 519560 474410
rect 519660 474310 519784 474410
rect 519884 474310 520008 474410
rect 520108 474310 520232 474410
rect 520332 474310 520456 474410
rect 520556 474310 520680 474410
rect 520780 474310 520904 474410
rect 521004 474310 521128 474410
rect 521228 474310 521352 474410
rect 521452 474310 521576 474410
rect 521676 474310 521800 474410
rect 521900 474310 522024 474410
rect 522124 474310 522248 474410
rect 522348 474310 522472 474410
rect 522572 474310 522696 474410
rect 522796 474310 522920 474410
rect 523020 474310 523144 474410
rect 523244 474310 523368 474410
rect 523468 474310 523592 474410
rect 523692 474310 523816 474410
rect 523916 474310 523940 474410
rect 530664 483236 537320 487356
rect 530664 478452 530760 483236
rect 536504 478452 537320 483236
rect 517260 474276 523940 474310
rect 527584 474280 528624 474336
rect 500364 474056 501404 474180
rect 511584 474212 511648 474276
rect 511712 474212 511776 474276
rect 511840 474212 511904 474276
rect 511968 474212 512032 474276
rect 512096 474212 512160 474276
rect 511584 474148 512160 474212
rect 527584 474180 527618 474280
rect 527718 474180 527842 474280
rect 527942 474180 528066 474280
rect 528166 474180 528290 474280
rect 528390 474180 528514 474280
rect 528614 474180 528624 474280
rect 500364 473956 500398 474056
rect 500498 473956 500622 474056
rect 500722 473956 500846 474056
rect 500946 473956 501070 474056
rect 501170 473956 501294 474056
rect 501394 473956 501404 474056
rect 500364 473832 501404 473956
rect 500364 473732 500398 473832
rect 500498 473732 500622 473832
rect 500722 473732 500846 473832
rect 500946 473732 501070 473832
rect 501170 473732 501294 473832
rect 501394 473732 501404 473832
rect 500364 473608 501404 473732
rect 500364 473508 500398 473608
rect 500498 473508 500622 473608
rect 500722 473508 500846 473608
rect 500946 473508 501070 473608
rect 501170 473508 501294 473608
rect 501394 473508 501404 473608
rect 500364 473384 501404 473508
rect 500364 473284 500398 473384
rect 500498 473284 500622 473384
rect 500722 473284 500846 473384
rect 500946 473284 501070 473384
rect 501170 473284 501294 473384
rect 501394 473284 501404 473384
rect 500364 473160 501404 473284
rect 500364 473060 500398 473160
rect 500498 473060 500622 473160
rect 500722 473060 500846 473160
rect 500946 473060 501070 473160
rect 501170 473060 501294 473160
rect 501394 473060 501404 473160
rect 500364 472936 501404 473060
rect 500364 472836 500398 472936
rect 500498 472836 500622 472936
rect 500722 472836 500846 472936
rect 500946 472836 501070 472936
rect 501170 472836 501294 472936
rect 501394 472836 501404 472936
rect 500364 472712 501404 472836
rect 500364 472612 500398 472712
rect 500498 472612 500622 472712
rect 500722 472612 500846 472712
rect 500946 472612 501070 472712
rect 501170 472612 501294 472712
rect 501394 472612 501404 472712
rect 500364 472488 501404 472612
rect 527584 474056 528624 474180
rect 527584 473956 527618 474056
rect 527718 473956 527842 474056
rect 527942 473956 528066 474056
rect 528166 473956 528290 474056
rect 528390 473956 528514 474056
rect 528614 473956 528624 474056
rect 527584 473832 528624 473956
rect 527584 473732 527618 473832
rect 527718 473732 527842 473832
rect 527942 473732 528066 473832
rect 528166 473732 528290 473832
rect 528390 473732 528514 473832
rect 528614 473732 528624 473832
rect 527584 473608 528624 473732
rect 527584 473508 527618 473608
rect 527718 473508 527842 473608
rect 527942 473508 528066 473608
rect 528166 473508 528290 473608
rect 528390 473508 528514 473608
rect 528614 473508 528624 473608
rect 527584 473384 528624 473508
rect 527584 473284 527618 473384
rect 527718 473284 527842 473384
rect 527942 473284 528066 473384
rect 528166 473284 528290 473384
rect 528390 473284 528514 473384
rect 528614 473284 528624 473384
rect 527584 473160 528624 473284
rect 527584 473060 527618 473160
rect 527718 473060 527842 473160
rect 527942 473060 528066 473160
rect 528166 473060 528290 473160
rect 528390 473060 528514 473160
rect 528614 473060 528624 473160
rect 527584 472936 528624 473060
rect 527584 472836 527618 472936
rect 527718 472836 527842 472936
rect 527942 472836 528066 472936
rect 528166 472836 528290 472936
rect 528390 472836 528514 472936
rect 528614 472836 528624 472936
rect 527584 472712 528624 472836
rect 527584 472612 527618 472712
rect 527718 472612 527842 472712
rect 527942 472612 528066 472712
rect 528166 472612 528290 472712
rect 528390 472612 528514 472712
rect 528614 472612 528624 472712
rect 500364 472388 500398 472488
rect 500498 472388 500622 472488
rect 500722 472388 500846 472488
rect 500946 472388 501070 472488
rect 501170 472388 501294 472488
rect 501394 472388 501404 472488
rect 518382 472513 526544 472530
rect 518382 472484 525651 472513
rect 500364 472264 501404 472388
rect 500364 472164 500398 472264
rect 500498 472164 500622 472264
rect 500722 472164 500846 472264
rect 500946 472164 501070 472264
rect 501170 472164 501294 472264
rect 501394 472164 501404 472264
rect 500364 472040 501404 472164
rect 500364 471940 500398 472040
rect 500498 471940 500622 472040
rect 500722 471940 500846 472040
rect 500946 471940 501070 472040
rect 501170 471940 501294 472040
rect 501394 471940 501404 472040
rect 500364 471816 501404 471940
rect 500364 471716 500398 471816
rect 500498 471716 500622 471816
rect 500722 471716 500846 471816
rect 500946 471716 501070 471816
rect 501170 471716 501294 471816
rect 501394 471716 501404 471816
rect 500364 471592 501404 471716
rect 500364 471492 500398 471592
rect 500498 471492 500622 471592
rect 500722 471492 500846 471592
rect 500946 471492 501070 471592
rect 501170 471492 501294 471592
rect 501394 471492 501404 471592
rect 500364 471368 501404 471492
rect 500364 471268 500398 471368
rect 500498 471268 500622 471368
rect 500722 471268 500846 471368
rect 500946 471268 501070 471368
rect 501170 471268 501294 471368
rect 501394 471268 501404 471368
rect 500364 471144 501404 471268
rect 500364 471044 500398 471144
rect 500498 471044 500622 471144
rect 500722 471044 500846 471144
rect 500946 471044 501070 471144
rect 501170 471044 501294 471144
rect 501394 471044 501404 471144
rect 500364 470920 501404 471044
rect 500364 470820 500398 470920
rect 500498 470820 500622 470920
rect 500722 470820 500846 470920
rect 500946 470820 501070 470920
rect 501170 470820 501294 470920
rect 501394 470820 501404 470920
rect 500364 470696 501404 470820
rect 500364 470596 500398 470696
rect 500498 470596 500622 470696
rect 500722 470596 500846 470696
rect 500946 470596 501070 470696
rect 501170 470596 501294 470696
rect 501394 470596 501404 470696
rect 500364 470472 501404 470596
rect 500364 470372 500398 470472
rect 500498 470372 500622 470472
rect 500722 470372 500846 470472
rect 500946 470372 501070 470472
rect 501170 470372 501294 470472
rect 501394 470372 501404 470472
rect 500364 470248 501404 470372
rect 500364 470148 500398 470248
rect 500498 470148 500622 470248
rect 500722 470148 500846 470248
rect 500946 470148 501070 470248
rect 501170 470148 501294 470248
rect 501394 470148 501404 470248
rect 500364 470024 501404 470148
rect 500364 469924 500398 470024
rect 500498 469924 500622 470024
rect 500722 469924 500846 470024
rect 500946 469924 501070 470024
rect 501170 469924 501294 470024
rect 501394 469924 501404 470024
rect 500364 469800 501404 469924
rect 500364 469700 500398 469800
rect 500498 469700 500622 469800
rect 500722 469700 500846 469800
rect 500946 469700 501070 469800
rect 501170 469700 501294 469800
rect 501394 469700 501404 469800
rect 500364 469576 501404 469700
rect 500364 469476 500398 469576
rect 500498 469476 500622 469576
rect 500722 469476 500846 469576
rect 500946 469476 501070 469576
rect 501170 469476 501294 469576
rect 501394 469476 501404 469576
rect 505787 469566 506071 469568
rect 500364 469352 501404 469476
rect 500364 469252 500398 469352
rect 500498 469252 500622 469352
rect 500722 469252 500846 469352
rect 500946 469252 501070 469352
rect 501170 469252 501294 469352
rect 501394 469252 501404 469352
rect 500364 469128 501404 469252
rect 500364 469028 500398 469128
rect 500498 469028 500622 469128
rect 500722 469028 500846 469128
rect 500946 469028 501070 469128
rect 501170 469028 501294 469128
rect 501394 469028 501404 469128
rect 500364 468904 501404 469028
rect 500364 468804 500398 468904
rect 500498 468804 500622 468904
rect 500722 468804 500846 468904
rect 500946 468804 501070 468904
rect 501170 468804 501294 468904
rect 501394 468804 501404 468904
rect 500364 468680 501404 468804
rect 500364 468580 500398 468680
rect 500498 468580 500622 468680
rect 500722 468580 500846 468680
rect 500946 468580 501070 468680
rect 501170 468580 501294 468680
rect 501394 468580 501404 468680
rect 500364 468456 501404 468580
rect 500364 468356 500398 468456
rect 500498 468356 500622 468456
rect 500722 468356 500846 468456
rect 500946 468356 501070 468456
rect 501170 468356 501294 468456
rect 501394 468356 501404 468456
rect 500364 468232 501404 468356
rect 500364 468132 500398 468232
rect 500498 468132 500622 468232
rect 500722 468132 500846 468232
rect 500946 468132 501070 468232
rect 501170 468132 501294 468232
rect 501394 468132 501404 468232
rect 500364 468008 501404 468132
rect 500364 467908 500398 468008
rect 500498 467908 500622 468008
rect 500722 467908 500846 468008
rect 500946 467908 501070 468008
rect 501170 467908 501294 468008
rect 501394 467908 501404 468008
rect 500364 467784 501404 467908
rect 500364 467684 500398 467784
rect 500498 467684 500622 467784
rect 500722 467684 500846 467784
rect 500946 467684 501070 467784
rect 501170 467684 501294 467784
rect 501394 467684 501404 467784
rect 500364 467680 501404 467684
rect 505786 468938 505789 469566
rect 506069 468938 511117 469566
rect 505786 468740 511117 468938
rect 505786 468700 517992 468740
rect 505786 468380 511332 468700
rect 511652 468380 512032 468700
rect 512352 468380 512732 468700
rect 513052 468380 513432 468700
rect 513752 468380 514132 468700
rect 514452 468380 514832 468700
rect 515152 468380 515532 468700
rect 515852 468380 516232 468700
rect 516552 468380 516932 468700
rect 517252 468380 517632 468700
rect 517952 468380 517992 468700
rect 505786 468340 517992 468380
rect 505786 468020 511124 468340
rect 511204 468225 511780 468241
rect 511204 468161 511220 468225
rect 511764 468161 511780 468225
rect 511204 468145 511780 468161
rect 511904 468225 512480 468241
rect 511904 468161 511920 468225
rect 512464 468161 512480 468225
rect 511904 468145 512480 468161
rect 512604 468225 513180 468241
rect 512604 468161 512620 468225
rect 513164 468161 513180 468225
rect 512604 468145 513180 468161
rect 513304 468225 513880 468241
rect 513304 468161 513320 468225
rect 513864 468161 513880 468225
rect 513304 468145 513880 468161
rect 514004 468225 514580 468241
rect 514004 468161 514020 468225
rect 514564 468161 514580 468225
rect 514004 468145 514580 468161
rect 514704 468225 515280 468241
rect 514704 468161 514720 468225
rect 515264 468161 515280 468225
rect 514704 468145 515280 468161
rect 515404 468225 515980 468241
rect 515404 468161 515420 468225
rect 515964 468161 515980 468225
rect 515404 468145 515980 468161
rect 516104 468225 516680 468241
rect 516104 468161 516120 468225
rect 516664 468161 516680 468225
rect 516104 468145 516680 468161
rect 516804 468225 517380 468241
rect 516804 468161 516820 468225
rect 517364 468161 517380 468225
rect 516804 468145 517380 468161
rect 517504 468225 518080 468241
rect 517504 468161 517520 468225
rect 518064 468161 518080 468225
rect 517504 468145 518080 468161
rect 505786 467981 517992 468020
rect 500393 467679 500503 467680
rect 500617 467679 500727 467680
rect 500841 467679 500951 467680
rect 501065 467679 501175 467680
rect 501289 467679 501399 467680
rect 505786 467661 511332 467981
rect 511652 467661 512032 467981
rect 512352 467661 512732 467981
rect 513052 467661 513432 467981
rect 513752 467661 514132 467981
rect 514452 467661 514832 467981
rect 515152 467661 515532 467981
rect 515852 467661 516232 467981
rect 516552 467661 516932 467981
rect 517252 467661 517632 467981
rect 517952 467661 517992 467981
rect 505786 467620 517992 467661
rect 505786 467300 511124 467620
rect 511204 467506 511780 467522
rect 511204 467442 511220 467506
rect 511764 467442 511780 467506
rect 511204 467426 511780 467442
rect 511904 467506 512480 467522
rect 511904 467442 511920 467506
rect 512464 467442 512480 467506
rect 511904 467426 512480 467442
rect 512604 467506 513180 467522
rect 512604 467442 512620 467506
rect 513164 467442 513180 467506
rect 512604 467426 513180 467442
rect 513304 467506 513880 467522
rect 513304 467442 513320 467506
rect 513864 467442 513880 467506
rect 513304 467426 513880 467442
rect 514004 467506 514580 467522
rect 514004 467442 514020 467506
rect 514564 467442 514580 467506
rect 514004 467426 514580 467442
rect 514704 467506 515280 467522
rect 514704 467442 514720 467506
rect 515264 467442 515280 467506
rect 514704 467426 515280 467442
rect 515404 467506 515980 467522
rect 515404 467442 515420 467506
rect 515964 467442 515980 467506
rect 515404 467426 515980 467442
rect 516104 467506 516680 467522
rect 516104 467442 516120 467506
rect 516664 467442 516680 467506
rect 516104 467426 516680 467442
rect 516804 467506 517380 467522
rect 516804 467442 516820 467506
rect 517364 467442 517380 467506
rect 516804 467426 517380 467442
rect 517504 467506 518080 467522
rect 517504 467442 517520 467506
rect 518064 467442 518080 467506
rect 517504 467426 518080 467442
rect 505786 467262 517992 467300
rect 505786 466942 511332 467262
rect 511652 466942 512032 467262
rect 512352 466942 512732 467262
rect 513052 466942 513432 467262
rect 513752 466942 514132 467262
rect 514452 466942 514832 467262
rect 515152 466942 515532 467262
rect 515852 466942 516232 467262
rect 516552 466942 516932 467262
rect 517252 466942 517632 467262
rect 517952 466942 517992 467262
rect 505786 466900 517992 466942
rect 505786 466580 511124 466900
rect 511204 466787 511780 466803
rect 511204 466723 511220 466787
rect 511764 466723 511780 466787
rect 511204 466707 511780 466723
rect 511904 466787 512480 466803
rect 511904 466723 511920 466787
rect 512464 466723 512480 466787
rect 511904 466707 512480 466723
rect 512604 466787 513180 466803
rect 512604 466723 512620 466787
rect 513164 466723 513180 466787
rect 512604 466707 513180 466723
rect 513304 466787 513880 466803
rect 513304 466723 513320 466787
rect 513864 466723 513880 466787
rect 513304 466707 513880 466723
rect 514004 466787 514580 466803
rect 514004 466723 514020 466787
rect 514564 466723 514580 466787
rect 514004 466707 514580 466723
rect 514704 466787 515280 466803
rect 514704 466723 514720 466787
rect 515264 466723 515280 466787
rect 514704 466707 515280 466723
rect 515404 466787 515980 466803
rect 515404 466723 515420 466787
rect 515964 466723 515980 466787
rect 515404 466707 515980 466723
rect 516104 466787 516680 466803
rect 516104 466723 516120 466787
rect 516664 466723 516680 466787
rect 516104 466707 516680 466723
rect 516804 466787 517380 466803
rect 516804 466723 516820 466787
rect 517364 466723 517380 466787
rect 516804 466707 517380 466723
rect 517504 466787 518080 466803
rect 517504 466723 517520 466787
rect 518064 466723 518080 466787
rect 517504 466707 518080 466723
rect 505786 466543 517992 466580
rect 505786 466223 511332 466543
rect 511652 466223 512032 466543
rect 512352 466223 512732 466543
rect 513052 466223 513432 466543
rect 513752 466223 514132 466543
rect 514452 466223 514832 466543
rect 515152 466223 515532 466543
rect 515852 466223 516232 466543
rect 516552 466223 516932 466543
rect 517252 466223 517632 466543
rect 517952 466223 517992 466543
rect 505786 466180 517992 466223
rect 505786 465860 511124 466180
rect 511204 466068 511780 466084
rect 511204 466004 511220 466068
rect 511764 466004 511780 466068
rect 511204 465988 511780 466004
rect 511904 466068 512480 466084
rect 511904 466004 511920 466068
rect 512464 466004 512480 466068
rect 511904 465988 512480 466004
rect 512604 466068 513180 466084
rect 512604 466004 512620 466068
rect 513164 466004 513180 466068
rect 512604 465988 513180 466004
rect 513304 466068 513880 466084
rect 513304 466004 513320 466068
rect 513864 466004 513880 466068
rect 513304 465988 513880 466004
rect 514004 466068 514580 466084
rect 514004 466004 514020 466068
rect 514564 466004 514580 466068
rect 514004 465988 514580 466004
rect 514704 466068 515280 466084
rect 514704 466004 514720 466068
rect 515264 466004 515280 466068
rect 514704 465988 515280 466004
rect 515404 466068 515980 466084
rect 515404 466004 515420 466068
rect 515964 466004 515980 466068
rect 515404 465988 515980 466004
rect 516104 466068 516680 466084
rect 516104 466004 516120 466068
rect 516664 466004 516680 466068
rect 516104 465988 516680 466004
rect 516804 466068 517380 466084
rect 516804 466004 516820 466068
rect 517364 466004 517380 466068
rect 516804 465988 517380 466004
rect 517504 466068 518080 466084
rect 517504 466004 517520 466068
rect 518064 466004 518080 466068
rect 517504 465988 518080 466004
rect 505786 465824 517992 465860
rect 505786 465504 511332 465824
rect 511652 465504 512032 465824
rect 512352 465504 512732 465824
rect 513052 465504 513432 465824
rect 513752 465504 514132 465824
rect 514452 465504 514832 465824
rect 515152 465504 515532 465824
rect 515852 465504 516232 465824
rect 516552 465504 516932 465824
rect 517252 465504 517632 465824
rect 517952 465504 517992 465824
rect 505786 465460 517992 465504
rect 505786 465140 511124 465460
rect 511204 465349 511780 465365
rect 511204 465285 511220 465349
rect 511764 465285 511780 465349
rect 511204 465269 511780 465285
rect 511904 465349 512480 465365
rect 511904 465285 511920 465349
rect 512464 465285 512480 465349
rect 511904 465269 512480 465285
rect 512604 465349 513180 465365
rect 512604 465285 512620 465349
rect 513164 465285 513180 465349
rect 512604 465269 513180 465285
rect 513304 465349 513880 465365
rect 513304 465285 513320 465349
rect 513864 465285 513880 465349
rect 513304 465269 513880 465285
rect 514004 465349 514580 465365
rect 514004 465285 514020 465349
rect 514564 465285 514580 465349
rect 514004 465269 514580 465285
rect 514704 465349 515280 465365
rect 514704 465285 514720 465349
rect 515264 465285 515280 465349
rect 514704 465269 515280 465285
rect 515404 465349 515980 465365
rect 515404 465285 515420 465349
rect 515964 465285 515980 465349
rect 515404 465269 515980 465285
rect 516104 465349 516680 465365
rect 516104 465285 516120 465349
rect 516664 465285 516680 465349
rect 516104 465269 516680 465285
rect 516804 465349 517380 465365
rect 516804 465285 516820 465349
rect 517364 465285 517380 465349
rect 516804 465269 517380 465285
rect 517504 465349 518080 465365
rect 517504 465285 517520 465349
rect 518064 465285 518080 465349
rect 517504 465269 518080 465285
rect 505786 465105 517992 465140
rect 505786 464785 511332 465105
rect 511652 464785 512032 465105
rect 512352 464785 512732 465105
rect 513052 464785 513432 465105
rect 513752 464785 514132 465105
rect 514452 464785 514832 465105
rect 515152 464785 515532 465105
rect 515852 464785 516232 465105
rect 516552 464785 516932 465105
rect 517252 464785 517632 465105
rect 517952 464785 517992 465105
rect 505786 464740 517992 464785
rect 505786 464420 511124 464740
rect 511204 464630 511780 464646
rect 511204 464566 511220 464630
rect 511764 464566 511780 464630
rect 511204 464550 511780 464566
rect 511904 464630 512480 464646
rect 511904 464566 511920 464630
rect 512464 464566 512480 464630
rect 511904 464550 512480 464566
rect 512604 464630 513180 464646
rect 512604 464566 512620 464630
rect 513164 464566 513180 464630
rect 512604 464550 513180 464566
rect 513304 464630 513880 464646
rect 513304 464566 513320 464630
rect 513864 464566 513880 464630
rect 513304 464550 513880 464566
rect 514004 464630 514580 464646
rect 514004 464566 514020 464630
rect 514564 464566 514580 464630
rect 514004 464550 514580 464566
rect 514704 464630 515280 464646
rect 514704 464566 514720 464630
rect 515264 464566 515280 464630
rect 514704 464550 515280 464566
rect 515404 464630 515980 464646
rect 515404 464566 515420 464630
rect 515964 464566 515980 464630
rect 515404 464550 515980 464566
rect 516104 464630 516680 464646
rect 516104 464566 516120 464630
rect 516664 464566 516680 464630
rect 516104 464550 516680 464566
rect 516804 464630 517380 464646
rect 516804 464566 516820 464630
rect 517364 464566 517380 464630
rect 516804 464550 517380 464566
rect 517504 464630 518080 464646
rect 517504 464566 517520 464630
rect 518064 464566 518080 464630
rect 517504 464550 518080 464566
rect 505786 464386 517992 464420
rect 505786 464066 511332 464386
rect 511652 464066 512032 464386
rect 512352 464066 512732 464386
rect 513052 464066 513432 464386
rect 513752 464066 514132 464386
rect 514452 464066 514832 464386
rect 515152 464066 515532 464386
rect 515852 464066 516232 464386
rect 516552 464066 516932 464386
rect 517252 464066 517632 464386
rect 517952 464066 517992 464386
rect 505786 464020 517992 464066
rect 490440 462236 497096 463452
rect 490440 457452 491256 462236
rect 497000 457452 497096 462236
rect 490440 456856 497096 457452
rect 500364 463810 501404 463866
rect 500364 463710 500398 463810
rect 500498 463710 500622 463810
rect 500722 463710 500846 463810
rect 500946 463710 501070 463810
rect 501170 463710 501294 463810
rect 501394 463710 501404 463810
rect 500364 463586 501404 463710
rect 500364 463486 500398 463586
rect 500498 463486 500622 463586
rect 500722 463486 500846 463586
rect 500946 463486 501070 463586
rect 501170 463486 501294 463586
rect 501394 463486 501404 463586
rect 500364 463362 501404 463486
rect 500364 463262 500398 463362
rect 500498 463262 500622 463362
rect 500722 463262 500846 463362
rect 500946 463262 501070 463362
rect 501170 463262 501294 463362
rect 501394 463262 501404 463362
rect 500364 463138 501404 463262
rect 500364 463038 500398 463138
rect 500498 463038 500622 463138
rect 500722 463038 500846 463138
rect 500946 463038 501070 463138
rect 501170 463038 501294 463138
rect 501394 463038 501404 463138
rect 500364 462914 501404 463038
rect 500364 462814 500398 462914
rect 500498 462814 500622 462914
rect 500722 462814 500846 462914
rect 500946 462814 501070 462914
rect 501170 462814 501294 462914
rect 501394 462814 501404 462914
rect 500364 462690 501404 462814
rect 500364 462590 500398 462690
rect 500498 462590 500622 462690
rect 500722 462590 500846 462690
rect 500946 462590 501070 462690
rect 501170 462590 501294 462690
rect 501394 462590 501404 462690
rect 500364 462466 501404 462590
rect 500364 462366 500398 462466
rect 500498 462366 500622 462466
rect 500722 462366 500846 462466
rect 500946 462366 501070 462466
rect 501170 462366 501294 462466
rect 501394 462366 501404 462466
rect 500364 462242 501404 462366
rect 500364 462142 500398 462242
rect 500498 462142 500622 462242
rect 500722 462142 500846 462242
rect 500946 462142 501070 462242
rect 501170 462142 501294 462242
rect 501394 462142 501404 462242
rect 500364 462018 501404 462142
rect 500364 461918 500398 462018
rect 500498 461918 500622 462018
rect 500722 461918 500846 462018
rect 500946 461918 501070 462018
rect 501170 461918 501294 462018
rect 501394 461918 501404 462018
rect 500364 461794 501404 461918
rect 500364 461694 500398 461794
rect 500498 461694 500622 461794
rect 500722 461694 500846 461794
rect 500946 461694 501070 461794
rect 501170 461694 501294 461794
rect 501394 461694 501404 461794
rect 500364 461570 501404 461694
rect 500364 461470 500398 461570
rect 500498 461470 500622 461570
rect 500722 461470 500846 461570
rect 500946 461470 501070 461570
rect 501170 461470 501294 461570
rect 501394 461470 501404 461570
rect 500364 461346 501404 461470
rect 500364 461246 500398 461346
rect 500498 461246 500622 461346
rect 500722 461246 500846 461346
rect 500946 461246 501070 461346
rect 501170 461246 501294 461346
rect 501394 461246 501404 461346
rect 500364 461122 501404 461246
rect 500364 461022 500398 461122
rect 500498 461022 500622 461122
rect 500722 461022 500846 461122
rect 500946 461022 501070 461122
rect 501170 461022 501294 461122
rect 501394 461022 501404 461122
rect 500364 460898 501404 461022
rect 500364 460798 500398 460898
rect 500498 460798 500622 460898
rect 500722 460798 500846 460898
rect 500946 460798 501070 460898
rect 501170 460798 501294 460898
rect 501394 460798 501404 460898
rect 500364 460674 501404 460798
rect 500364 460574 500398 460674
rect 500498 460574 500622 460674
rect 500722 460574 500846 460674
rect 500946 460574 501070 460674
rect 501170 460574 501294 460674
rect 501394 460574 501404 460674
rect 500364 460450 501404 460574
rect 500364 460350 500398 460450
rect 500498 460350 500622 460450
rect 500722 460350 500846 460450
rect 500946 460350 501070 460450
rect 501170 460350 501294 460450
rect 501394 460350 501404 460450
rect 505786 463700 511124 464020
rect 511204 463911 511780 463927
rect 511204 463847 511220 463911
rect 511764 463847 511780 463911
rect 511204 463831 511780 463847
rect 511904 463911 512480 463927
rect 511904 463847 511920 463911
rect 512464 463847 512480 463911
rect 511904 463831 512480 463847
rect 512604 463911 513180 463927
rect 512604 463847 512620 463911
rect 513164 463847 513180 463911
rect 512604 463831 513180 463847
rect 513304 463911 513880 463927
rect 513304 463847 513320 463911
rect 513864 463847 513880 463911
rect 513304 463831 513880 463847
rect 514004 463911 514580 463927
rect 514004 463847 514020 463911
rect 514564 463847 514580 463911
rect 514004 463831 514580 463847
rect 514704 463911 515280 463927
rect 514704 463847 514720 463911
rect 515264 463847 515280 463911
rect 514704 463831 515280 463847
rect 515404 463911 515980 463927
rect 515404 463847 515420 463911
rect 515964 463847 515980 463911
rect 515404 463831 515980 463847
rect 516104 463911 516680 463927
rect 516104 463847 516120 463911
rect 516664 463847 516680 463911
rect 516104 463831 516680 463847
rect 516804 463911 517380 463927
rect 516804 463847 516820 463911
rect 517364 463847 517380 463911
rect 516804 463831 517380 463847
rect 517504 463911 518080 463927
rect 517504 463847 517520 463911
rect 518064 463847 518080 463911
rect 517504 463831 518080 463847
rect 505786 463667 517992 463700
rect 505786 463347 511332 463667
rect 511652 463347 512032 463667
rect 512352 463347 512732 463667
rect 513052 463347 513432 463667
rect 513752 463347 514132 463667
rect 514452 463347 514832 463667
rect 515152 463347 515532 463667
rect 515852 463347 516232 463667
rect 516552 463347 516932 463667
rect 517252 463347 517632 463667
rect 517952 463347 517992 463667
rect 505786 463300 517992 463347
rect 505786 462980 511124 463300
rect 511204 463192 511780 463208
rect 511204 463128 511220 463192
rect 511764 463128 511780 463192
rect 511204 463112 511780 463128
rect 511904 463192 512480 463208
rect 511904 463128 511920 463192
rect 512464 463128 512480 463192
rect 511904 463112 512480 463128
rect 512604 463192 513180 463208
rect 512604 463128 512620 463192
rect 513164 463128 513180 463192
rect 512604 463112 513180 463128
rect 513304 463192 513880 463208
rect 513304 463128 513320 463192
rect 513864 463128 513880 463192
rect 513304 463112 513880 463128
rect 514004 463192 514580 463208
rect 514004 463128 514020 463192
rect 514564 463128 514580 463192
rect 514004 463112 514580 463128
rect 514704 463192 515280 463208
rect 514704 463128 514720 463192
rect 515264 463128 515280 463192
rect 514704 463112 515280 463128
rect 515404 463192 515980 463208
rect 515404 463128 515420 463192
rect 515964 463128 515980 463192
rect 515404 463112 515980 463128
rect 516104 463192 516680 463208
rect 516104 463128 516120 463192
rect 516664 463128 516680 463192
rect 516104 463112 516680 463128
rect 516804 463192 517380 463208
rect 516804 463128 516820 463192
rect 517364 463128 517380 463192
rect 516804 463112 517380 463128
rect 517504 463192 518080 463208
rect 517504 463128 517520 463192
rect 518064 463128 518080 463192
rect 517504 463112 518080 463128
rect 505786 462948 517992 462980
rect 505786 462628 511332 462948
rect 511652 462628 512032 462948
rect 512352 462628 512732 462948
rect 513052 462628 513432 462948
rect 513752 462628 514132 462948
rect 514452 462628 514832 462948
rect 515152 462628 515532 462948
rect 515852 462628 516232 462948
rect 516552 462628 516932 462948
rect 517252 462628 517632 462948
rect 517952 462628 517992 462948
rect 505786 462580 517992 462628
rect 505786 462260 511124 462580
rect 511204 462473 511780 462489
rect 511204 462409 511220 462473
rect 511764 462409 511780 462473
rect 511204 462393 511780 462409
rect 511904 462473 512480 462489
rect 511904 462409 511920 462473
rect 512464 462409 512480 462473
rect 511904 462393 512480 462409
rect 512604 462473 513180 462489
rect 512604 462409 512620 462473
rect 513164 462409 513180 462473
rect 512604 462393 513180 462409
rect 513304 462473 513880 462489
rect 513304 462409 513320 462473
rect 513864 462409 513880 462473
rect 513304 462393 513880 462409
rect 514004 462473 514580 462489
rect 514004 462409 514020 462473
rect 514564 462409 514580 462473
rect 514004 462393 514580 462409
rect 514704 462473 515280 462489
rect 514704 462409 514720 462473
rect 515264 462409 515280 462473
rect 514704 462393 515280 462409
rect 515404 462473 515980 462489
rect 515404 462409 515420 462473
rect 515964 462409 515980 462473
rect 515404 462393 515980 462409
rect 516104 462473 516680 462489
rect 516104 462409 516120 462473
rect 516664 462409 516680 462473
rect 516104 462393 516680 462409
rect 516804 462473 517380 462489
rect 516804 462409 516820 462473
rect 517364 462409 517380 462473
rect 516804 462393 517380 462409
rect 517504 462473 518080 462489
rect 517504 462409 517520 462473
rect 518064 462409 518080 462473
rect 517504 462393 518080 462409
rect 517592 462260 517992 462269
rect 505786 462229 517992 462260
rect 505786 461909 511332 462229
rect 511652 461909 512032 462229
rect 512352 461909 512732 462229
rect 513052 461909 513432 462229
rect 513752 461909 514132 462229
rect 514452 461909 514832 462229
rect 515152 461909 515532 462229
rect 515852 461909 516232 462229
rect 516552 461909 516932 462229
rect 517252 461909 517632 462229
rect 517952 461909 517992 462229
rect 505786 461860 517992 461909
rect 505786 461840 511132 461860
rect 505786 461075 511117 461840
rect 511204 461754 511780 461770
rect 511204 461690 511220 461754
rect 511764 461690 511780 461754
rect 511204 461674 511780 461690
rect 511904 461754 512480 461770
rect 511904 461690 511920 461754
rect 512464 461690 512480 461754
rect 511904 461674 512480 461690
rect 512604 461754 513180 461770
rect 512604 461690 512620 461754
rect 513164 461690 513180 461754
rect 512604 461674 513180 461690
rect 513304 461754 513880 461770
rect 513304 461690 513320 461754
rect 513864 461690 513880 461754
rect 513304 461674 513880 461690
rect 514004 461754 514580 461770
rect 514004 461690 514020 461754
rect 514564 461690 514580 461754
rect 514004 461674 514580 461690
rect 514704 461754 515280 461770
rect 514704 461690 514720 461754
rect 515264 461690 515280 461754
rect 514704 461674 515280 461690
rect 515404 461754 515980 461770
rect 515404 461690 515420 461754
rect 515964 461690 515980 461754
rect 515404 461674 515980 461690
rect 516104 461754 516680 461770
rect 516104 461690 516120 461754
rect 516664 461690 516680 461754
rect 516104 461674 516680 461690
rect 516804 461754 517380 461770
rect 516804 461690 516820 461754
rect 517364 461690 517380 461754
rect 516804 461674 517380 461690
rect 517504 461754 518080 461770
rect 517504 461690 517520 461754
rect 518064 461690 518080 461754
rect 517504 461674 518080 461690
rect 518376 461239 525651 472484
rect 526507 461239 526544 472513
rect 527584 472488 528624 472612
rect 527584 472388 527618 472488
rect 527718 472388 527842 472488
rect 527942 472388 528066 472488
rect 528166 472388 528290 472488
rect 528390 472388 528514 472488
rect 528614 472388 528624 472488
rect 527584 472264 528624 472388
rect 527584 472164 527618 472264
rect 527718 472164 527842 472264
rect 527942 472164 528066 472264
rect 528166 472164 528290 472264
rect 528390 472164 528514 472264
rect 528614 472164 528624 472264
rect 527584 472040 528624 472164
rect 527584 471940 527618 472040
rect 527718 471940 527842 472040
rect 527942 471940 528066 472040
rect 528166 471940 528290 472040
rect 528390 471940 528514 472040
rect 528614 471940 528624 472040
rect 527584 471816 528624 471940
rect 527584 471716 527618 471816
rect 527718 471716 527842 471816
rect 527942 471716 528066 471816
rect 528166 471716 528290 471816
rect 528390 471716 528514 471816
rect 528614 471716 528624 471816
rect 527584 471592 528624 471716
rect 527584 471492 527618 471592
rect 527718 471492 527842 471592
rect 527942 471492 528066 471592
rect 528166 471492 528290 471592
rect 528390 471492 528514 471592
rect 528614 471492 528624 471592
rect 527584 471368 528624 471492
rect 527584 471268 527618 471368
rect 527718 471268 527842 471368
rect 527942 471268 528066 471368
rect 528166 471268 528290 471368
rect 528390 471268 528514 471368
rect 528614 471268 528624 471368
rect 527584 471144 528624 471268
rect 527584 471044 527618 471144
rect 527718 471044 527842 471144
rect 527942 471044 528066 471144
rect 528166 471044 528290 471144
rect 528390 471044 528514 471144
rect 528614 471044 528624 471144
rect 527584 470920 528624 471044
rect 527584 470820 527618 470920
rect 527718 470820 527842 470920
rect 527942 470820 528066 470920
rect 528166 470820 528290 470920
rect 528390 470820 528514 470920
rect 528614 470820 528624 470920
rect 527584 470696 528624 470820
rect 527584 470596 527618 470696
rect 527718 470596 527842 470696
rect 527942 470596 528066 470696
rect 528166 470596 528290 470696
rect 528390 470596 528514 470696
rect 528614 470596 528624 470696
rect 527584 470472 528624 470596
rect 527584 470372 527618 470472
rect 527718 470372 527842 470472
rect 527942 470372 528066 470472
rect 528166 470372 528290 470472
rect 528390 470372 528514 470472
rect 528614 470372 528624 470472
rect 527584 470248 528624 470372
rect 527584 470148 527618 470248
rect 527718 470148 527842 470248
rect 527942 470148 528066 470248
rect 528166 470148 528290 470248
rect 528390 470148 528514 470248
rect 528614 470148 528624 470248
rect 527584 470024 528624 470148
rect 527584 469924 527618 470024
rect 527718 469924 527842 470024
rect 527942 469924 528066 470024
rect 528166 469924 528290 470024
rect 528390 469924 528514 470024
rect 528614 469924 528624 470024
rect 527584 469800 528624 469924
rect 527584 469700 527618 469800
rect 527718 469700 527842 469800
rect 527942 469700 528066 469800
rect 528166 469700 528290 469800
rect 528390 469700 528514 469800
rect 528614 469700 528624 469800
rect 527584 469576 528624 469700
rect 527584 469476 527618 469576
rect 527718 469476 527842 469576
rect 527942 469476 528066 469576
rect 528166 469476 528290 469576
rect 528390 469476 528514 469576
rect 528614 469476 528624 469576
rect 527584 469352 528624 469476
rect 527584 469252 527618 469352
rect 527718 469252 527842 469352
rect 527942 469252 528066 469352
rect 528166 469252 528290 469352
rect 528390 469252 528514 469352
rect 528614 469252 528624 469352
rect 527584 469128 528624 469252
rect 527584 469028 527618 469128
rect 527718 469028 527842 469128
rect 527942 469028 528066 469128
rect 528166 469028 528290 469128
rect 528390 469028 528514 469128
rect 528614 469028 528624 469128
rect 527584 468904 528624 469028
rect 527584 468804 527618 468904
rect 527718 468804 527842 468904
rect 527942 468804 528066 468904
rect 528166 468804 528290 468904
rect 528390 468804 528514 468904
rect 528614 468804 528624 468904
rect 527584 468680 528624 468804
rect 527584 468580 527618 468680
rect 527718 468580 527842 468680
rect 527942 468580 528066 468680
rect 528166 468580 528290 468680
rect 528390 468580 528514 468680
rect 528614 468580 528624 468680
rect 527584 468456 528624 468580
rect 527584 468356 527618 468456
rect 527718 468356 527842 468456
rect 527942 468356 528066 468456
rect 528166 468356 528290 468456
rect 528390 468356 528514 468456
rect 528614 468356 528624 468456
rect 527584 468232 528624 468356
rect 527584 468132 527618 468232
rect 527718 468132 527842 468232
rect 527942 468132 528066 468232
rect 528166 468132 528290 468232
rect 528390 468132 528514 468232
rect 528614 468132 528624 468232
rect 527584 468008 528624 468132
rect 527584 467908 527618 468008
rect 527718 467908 527842 468008
rect 527942 467908 528066 468008
rect 528166 467908 528290 468008
rect 528390 467908 528514 468008
rect 528614 467908 528624 468008
rect 527584 467784 528624 467908
rect 527584 467684 527618 467784
rect 527718 467684 527842 467784
rect 527942 467684 528066 467784
rect 528166 467684 528290 467784
rect 528390 467684 528514 467784
rect 528614 467684 528624 467784
rect 527584 467680 528624 467684
rect 530664 474236 537320 478452
rect 572536 484036 577492 484272
rect 572536 477664 572772 484036
rect 573008 477664 573244 484036
rect 573480 477664 573716 484036
rect 573952 477664 574188 484036
rect 574424 477664 574660 484036
rect 574896 477664 575132 484036
rect 575368 477664 575604 484036
rect 575840 477664 576076 484036
rect 576312 477664 576548 484036
rect 576784 477664 577020 484036
rect 577256 477664 577492 484036
rect 530664 469452 530760 474236
rect 536504 469452 537320 474236
rect 530664 468236 537320 469452
rect 527613 467679 527723 467680
rect 527837 467679 527947 467680
rect 528061 467679 528171 467680
rect 528285 467679 528395 467680
rect 528509 467679 528619 467680
rect 518376 461204 526544 461239
rect 527584 463810 528624 463866
rect 527584 463710 527618 463810
rect 527718 463710 527842 463810
rect 527942 463710 528066 463810
rect 528166 463710 528290 463810
rect 528390 463710 528514 463810
rect 528614 463710 528624 463810
rect 527584 463586 528624 463710
rect 527584 463486 527618 463586
rect 527718 463486 527842 463586
rect 527942 463486 528066 463586
rect 528166 463486 528290 463586
rect 528390 463486 528514 463586
rect 528614 463486 528624 463586
rect 527584 463362 528624 463486
rect 527584 463262 527618 463362
rect 527718 463262 527842 463362
rect 527942 463262 528066 463362
rect 528166 463262 528290 463362
rect 528390 463262 528514 463362
rect 528614 463262 528624 463362
rect 527584 463138 528624 463262
rect 527584 463038 527618 463138
rect 527718 463038 527842 463138
rect 527942 463038 528066 463138
rect 528166 463038 528290 463138
rect 528390 463038 528514 463138
rect 528614 463038 528624 463138
rect 527584 462914 528624 463038
rect 527584 462814 527618 462914
rect 527718 462814 527842 462914
rect 527942 462814 528066 462914
rect 528166 462814 528290 462914
rect 528390 462814 528514 462914
rect 528614 462814 528624 462914
rect 527584 462690 528624 462814
rect 527584 462590 527618 462690
rect 527718 462590 527842 462690
rect 527942 462590 528066 462690
rect 528166 462590 528290 462690
rect 528390 462590 528514 462690
rect 528614 462590 528624 462690
rect 527584 462466 528624 462590
rect 527584 462366 527618 462466
rect 527718 462366 527842 462466
rect 527942 462366 528066 462466
rect 528166 462366 528290 462466
rect 528390 462366 528514 462466
rect 528614 462366 528624 462466
rect 527584 462242 528624 462366
rect 527584 462142 527618 462242
rect 527718 462142 527842 462242
rect 527942 462142 528066 462242
rect 528166 462142 528290 462242
rect 528390 462142 528514 462242
rect 528614 462142 528624 462242
rect 527584 462018 528624 462142
rect 527584 461918 527618 462018
rect 527718 461918 527842 462018
rect 527942 461918 528066 462018
rect 528166 461918 528290 462018
rect 528390 461918 528514 462018
rect 528614 461918 528624 462018
rect 527584 461794 528624 461918
rect 527584 461694 527618 461794
rect 527718 461694 527842 461794
rect 527942 461694 528066 461794
rect 528166 461694 528290 461794
rect 528390 461694 528514 461794
rect 528614 461694 528624 461794
rect 527584 461570 528624 461694
rect 527584 461470 527618 461570
rect 527718 461470 527842 461570
rect 527942 461470 528066 461570
rect 528166 461470 528290 461570
rect 528390 461470 528514 461570
rect 528614 461470 528624 461570
rect 527584 461346 528624 461470
rect 527584 461246 527618 461346
rect 527718 461246 527842 461346
rect 527942 461246 528066 461346
rect 528166 461246 528290 461346
rect 528390 461246 528514 461346
rect 528614 461246 528624 461346
rect 505786 460447 505789 461075
rect 506069 460447 511117 461075
rect 505786 460434 511117 460447
rect 527584 461122 528624 461246
rect 527584 461022 527618 461122
rect 527718 461022 527842 461122
rect 527942 461022 528066 461122
rect 528166 461022 528290 461122
rect 528390 461022 528514 461122
rect 528614 461022 528624 461122
rect 527584 460898 528624 461022
rect 527584 460798 527618 460898
rect 527718 460798 527842 460898
rect 527942 460798 528066 460898
rect 528166 460798 528290 460898
rect 528390 460798 528514 460898
rect 528614 460798 528624 460898
rect 527584 460674 528624 460798
rect 527584 460574 527618 460674
rect 527718 460574 527842 460674
rect 527942 460574 528066 460674
rect 528166 460574 528290 460674
rect 528390 460574 528514 460674
rect 528614 460574 528624 460674
rect 527584 460450 528624 460574
rect 500364 460226 501404 460350
rect 500364 460126 500398 460226
rect 500498 460126 500622 460226
rect 500722 460126 500846 460226
rect 500946 460126 501070 460226
rect 501170 460126 501294 460226
rect 501394 460126 501404 460226
rect 527584 460350 527618 460450
rect 527718 460350 527842 460450
rect 527942 460350 528066 460450
rect 528166 460350 528290 460450
rect 528390 460350 528514 460450
rect 528614 460350 528624 460450
rect 527584 460226 528624 460350
rect 500364 460002 501404 460126
rect 500364 459902 500398 460002
rect 500498 459902 500622 460002
rect 500722 459902 500846 460002
rect 500946 459902 501070 460002
rect 501170 459902 501294 460002
rect 501394 459902 501404 460002
rect 500364 459778 501404 459902
rect 500364 459678 500398 459778
rect 500498 459678 500622 459778
rect 500722 459678 500846 459778
rect 500946 459678 501070 459778
rect 501170 459678 501294 459778
rect 501394 459678 501404 459778
rect 500364 459554 501404 459678
rect 500364 459454 500398 459554
rect 500498 459454 500622 459554
rect 500722 459454 500846 459554
rect 500946 459454 501070 459554
rect 501170 459454 501294 459554
rect 501394 459454 501404 459554
rect 500364 459330 501404 459454
rect 500364 459230 500398 459330
rect 500498 459230 500622 459330
rect 500722 459230 500846 459330
rect 500946 459230 501070 459330
rect 501170 459230 501294 459330
rect 501394 459230 501404 459330
rect 500364 459106 501404 459230
rect 500364 459006 500398 459106
rect 500498 459006 500622 459106
rect 500722 459006 500846 459106
rect 500946 459006 501070 459106
rect 501170 459006 501294 459106
rect 501394 459006 501404 459106
rect 500364 458882 501404 459006
rect 500364 458782 500398 458882
rect 500498 458782 500622 458882
rect 500722 458782 500846 458882
rect 500946 458782 501070 458882
rect 501170 458782 501294 458882
rect 501394 458782 501404 458882
rect 500364 458658 501404 458782
rect 500364 458558 500398 458658
rect 500498 458558 500622 458658
rect 500722 458558 500846 458658
rect 500946 458558 501070 458658
rect 501170 458558 501294 458658
rect 501394 458558 501404 458658
rect 500364 458434 501404 458558
rect 500364 458334 500398 458434
rect 500498 458334 500622 458434
rect 500722 458334 500846 458434
rect 500946 458334 501070 458434
rect 501170 458334 501294 458434
rect 501394 458334 501404 458434
rect 500364 458210 501404 458334
rect 500364 458110 500398 458210
rect 500498 458110 500622 458210
rect 500722 458110 500846 458210
rect 500946 458110 501070 458210
rect 501170 458110 501294 458210
rect 501394 458110 501404 458210
rect 500364 457986 501404 458110
rect 500364 457886 500398 457986
rect 500498 457886 500622 457986
rect 500722 457886 500846 457986
rect 500946 457886 501070 457986
rect 501170 457886 501294 457986
rect 501394 457886 501404 457986
rect 500364 457762 501404 457886
rect 500364 457662 500398 457762
rect 500498 457662 500622 457762
rect 500722 457662 500846 457762
rect 500946 457662 501070 457762
rect 501170 457662 501294 457762
rect 501394 457662 501404 457762
rect 500364 457538 501404 457662
rect 500364 457438 500398 457538
rect 500498 457438 500622 457538
rect 500722 457438 500846 457538
rect 500946 457438 501070 457538
rect 501170 457438 501294 457538
rect 501394 457438 501404 457538
rect 500364 457314 501404 457438
rect 500364 457214 500398 457314
rect 500498 457214 500622 457314
rect 500722 457214 500846 457314
rect 500946 457214 501070 457314
rect 501170 457214 501294 457314
rect 501394 457214 501404 457314
rect 500364 457210 501404 457214
rect 512233 460198 513207 460199
rect 500393 457209 500503 457210
rect 500617 457209 500727 457210
rect 500841 457209 500951 457210
rect 501065 457209 501175 457210
rect 501289 457209 501399 457210
rect 477060 450892 477500 455676
rect 483244 450892 483726 455676
rect 477060 447676 483726 450892
rect 477060 442892 477500 447676
rect 483244 442892 483726 447676
rect 477060 378072 483726 442892
rect 490464 436676 497126 456856
rect 512233 439888 512234 460198
rect 513206 439888 513207 460198
rect 527584 460126 527618 460226
rect 527718 460126 527842 460226
rect 527942 460126 528066 460226
rect 528166 460126 528290 460226
rect 528390 460126 528514 460226
rect 528614 460126 528624 460226
rect 527584 460002 528624 460126
rect 527584 459902 527618 460002
rect 527718 459902 527842 460002
rect 527942 459902 528066 460002
rect 528166 459902 528290 460002
rect 528390 459902 528514 460002
rect 528614 459902 528624 460002
rect 527584 459778 528624 459902
rect 527584 459678 527618 459778
rect 527718 459678 527842 459778
rect 527942 459678 528066 459778
rect 528166 459678 528290 459778
rect 528390 459678 528514 459778
rect 528614 459678 528624 459778
rect 527584 459554 528624 459678
rect 527584 459454 527618 459554
rect 527718 459454 527842 459554
rect 527942 459454 528066 459554
rect 528166 459454 528290 459554
rect 528390 459454 528514 459554
rect 528614 459454 528624 459554
rect 527584 459330 528624 459454
rect 527584 459230 527618 459330
rect 527718 459230 527842 459330
rect 527942 459230 528066 459330
rect 528166 459230 528290 459330
rect 528390 459230 528514 459330
rect 528614 459230 528624 459330
rect 527584 459106 528624 459230
rect 527584 459006 527618 459106
rect 527718 459006 527842 459106
rect 527942 459006 528066 459106
rect 528166 459006 528290 459106
rect 528390 459006 528514 459106
rect 528614 459006 528624 459106
rect 527584 458882 528624 459006
rect 527584 458782 527618 458882
rect 527718 458782 527842 458882
rect 527942 458782 528066 458882
rect 528166 458782 528290 458882
rect 528390 458782 528514 458882
rect 528614 458782 528624 458882
rect 527584 458658 528624 458782
rect 527584 458558 527618 458658
rect 527718 458558 527842 458658
rect 527942 458558 528066 458658
rect 528166 458558 528290 458658
rect 528390 458558 528514 458658
rect 528614 458558 528624 458658
rect 527584 458434 528624 458558
rect 527584 458334 527618 458434
rect 527718 458334 527842 458434
rect 527942 458334 528066 458434
rect 528166 458334 528290 458434
rect 528390 458334 528514 458434
rect 528614 458334 528624 458434
rect 527584 458210 528624 458334
rect 527584 458110 527618 458210
rect 527718 458110 527842 458210
rect 527942 458110 528066 458210
rect 528166 458110 528290 458210
rect 528390 458110 528514 458210
rect 528614 458110 528624 458210
rect 527584 457986 528624 458110
rect 527584 457886 527618 457986
rect 527718 457886 527842 457986
rect 527942 457886 528066 457986
rect 528166 457886 528290 457986
rect 528390 457886 528514 457986
rect 528614 457886 528624 457986
rect 527584 457762 528624 457886
rect 527584 457662 527618 457762
rect 527718 457662 527842 457762
rect 527942 457662 528066 457762
rect 528166 457662 528290 457762
rect 528390 457662 528514 457762
rect 528614 457662 528624 457762
rect 527584 457538 528624 457662
rect 527584 457438 527618 457538
rect 527718 457438 527842 457538
rect 527942 457438 528066 457538
rect 528166 457438 528290 457538
rect 528390 457438 528514 457538
rect 528614 457438 528624 457538
rect 527584 457314 528624 457438
rect 527584 457214 527618 457314
rect 527718 457214 527842 457314
rect 527942 457214 528066 457314
rect 528166 457214 528290 457314
rect 528390 457214 528514 457314
rect 528614 457214 528624 457314
rect 527584 457210 528624 457214
rect 530664 463452 530760 468236
rect 536504 463452 537320 468236
rect 530664 462236 537320 463452
rect 530664 457452 530760 462236
rect 536504 457452 537320 462236
rect 527613 457209 527723 457210
rect 527837 457209 527947 457210
rect 528061 457209 528171 457210
rect 528285 457209 528395 457210
rect 528509 457209 528619 457210
rect 513719 453756 513921 453757
rect 513719 453556 513720 453756
rect 513920 453556 513921 453756
rect 513719 453555 513921 453556
rect 514153 453756 514355 453757
rect 514153 453556 514154 453756
rect 514354 453556 514355 453756
rect 514153 453555 514355 453556
rect 514587 453756 514789 453757
rect 514587 453556 514588 453756
rect 514788 453556 514789 453756
rect 514587 453555 514789 453556
rect 513719 453322 513921 453323
rect 513719 453122 513720 453322
rect 513920 453122 513921 453322
rect 513719 453121 513921 453122
rect 514153 453322 514355 453323
rect 514153 453122 514154 453322
rect 514354 453122 514355 453322
rect 514153 453121 514355 453122
rect 514587 453322 514789 453323
rect 514587 453122 514588 453322
rect 514788 453122 514789 453322
rect 514587 453121 514789 453122
rect 513719 452888 513921 452889
rect 513719 452688 513720 452888
rect 513920 452688 513921 452888
rect 513719 452687 513921 452688
rect 514153 452888 514355 452889
rect 514153 452688 514154 452888
rect 514354 452688 514355 452888
rect 514153 452687 514355 452688
rect 514587 452888 514789 452889
rect 514587 452688 514588 452888
rect 514788 452688 514789 452888
rect 514587 452687 514789 452688
rect 513719 452454 513921 452455
rect 513719 452254 513720 452454
rect 513920 452254 513921 452454
rect 513719 452253 513921 452254
rect 514153 452454 514355 452455
rect 514153 452254 514154 452454
rect 514354 452254 514355 452454
rect 514153 452253 514355 452254
rect 514587 452454 514789 452455
rect 514587 452254 514588 452454
rect 514788 452254 514789 452454
rect 514587 452253 514789 452254
rect 513719 452020 513921 452021
rect 513719 451820 513720 452020
rect 513920 451820 513921 452020
rect 513719 451819 513921 451820
rect 514153 452020 514355 452021
rect 514153 451820 514154 452020
rect 514354 451820 514355 452020
rect 514153 451819 514355 451820
rect 514587 452020 514789 452021
rect 514587 451820 514588 452020
rect 514788 451820 514789 452020
rect 514587 451819 514789 451820
rect 513719 451586 513921 451587
rect 513719 451386 513720 451586
rect 513920 451386 513921 451586
rect 513719 451385 513921 451386
rect 514153 451586 514355 451587
rect 514153 451386 514154 451586
rect 514354 451386 514355 451586
rect 514153 451385 514355 451386
rect 514587 451586 514789 451587
rect 514587 451386 514588 451586
rect 514788 451386 514789 451586
rect 514587 451385 514789 451386
rect 513719 451152 513921 451153
rect 513719 450952 513720 451152
rect 513920 450952 513921 451152
rect 513719 450951 513921 450952
rect 514153 451152 514355 451153
rect 514153 450952 514154 451152
rect 514354 450952 514355 451152
rect 514153 450951 514355 450952
rect 514587 451152 514789 451153
rect 514587 450952 514588 451152
rect 514788 450952 514789 451152
rect 514587 450951 514789 450952
rect 513719 450718 513921 450719
rect 513719 450518 513720 450718
rect 513920 450518 513921 450718
rect 513719 450517 513921 450518
rect 514153 450718 514355 450719
rect 514153 450518 514154 450718
rect 514354 450518 514355 450718
rect 514153 450517 514355 450518
rect 514587 450718 514789 450719
rect 514587 450518 514588 450718
rect 514788 450518 514789 450718
rect 514587 450517 514789 450518
rect 513719 450284 513921 450285
rect 513719 450084 513720 450284
rect 513920 450084 513921 450284
rect 513719 450083 513921 450084
rect 514153 450284 514355 450285
rect 514153 450084 514154 450284
rect 514354 450084 514355 450284
rect 514153 450083 514355 450084
rect 514587 450284 514789 450285
rect 514587 450084 514588 450284
rect 514788 450084 514789 450284
rect 514587 450083 514789 450084
rect 513719 449850 513921 449851
rect 513719 449650 513720 449850
rect 513920 449650 513921 449850
rect 513719 449649 513921 449650
rect 514153 449850 514355 449851
rect 514153 449650 514154 449850
rect 514354 449650 514355 449850
rect 514153 449649 514355 449650
rect 514587 449850 514789 449851
rect 514587 449650 514588 449850
rect 514788 449650 514789 449850
rect 514587 449649 514789 449650
rect 513719 449416 513921 449417
rect 513719 449216 513720 449416
rect 513920 449216 513921 449416
rect 513719 449215 513921 449216
rect 514153 449416 514355 449417
rect 514153 449216 514154 449416
rect 514354 449216 514355 449416
rect 514153 449215 514355 449216
rect 514587 449416 514789 449417
rect 514587 449216 514588 449416
rect 514788 449216 514789 449416
rect 514587 449215 514789 449216
rect 514587 449016 514789 449017
rect 514587 448816 514588 449016
rect 514788 448816 514789 449016
rect 514587 448815 514789 448816
rect 514587 448616 514789 448617
rect 514587 448416 514588 448616
rect 514788 448416 514789 448616
rect 514587 448415 514789 448416
rect 514587 448216 514789 448217
rect 514587 448016 514588 448216
rect 514788 448016 514789 448216
rect 514587 448015 514789 448016
rect 514587 447816 514789 447817
rect 514587 447616 514588 447816
rect 514788 447616 514789 447816
rect 514587 447615 514789 447616
rect 514587 447416 514789 447417
rect 514587 447216 514588 447416
rect 514788 447216 514789 447416
rect 514587 447215 514789 447216
rect 514587 447016 514789 447017
rect 514587 446816 514588 447016
rect 514788 446816 514789 447016
rect 514587 446815 514789 446816
rect 514587 446616 514789 446617
rect 514587 446416 514588 446616
rect 514788 446416 514789 446616
rect 514587 446415 514789 446416
rect 514587 446216 514789 446217
rect 514587 446016 514588 446216
rect 514788 446016 514789 446216
rect 514587 446015 514789 446016
rect 514587 445816 514789 445817
rect 514587 445616 514588 445816
rect 514788 445616 514789 445816
rect 514587 445615 514789 445616
rect 514587 444216 514789 444217
rect 514587 444016 514588 444216
rect 514788 444016 514789 444216
rect 514587 444015 514789 444016
rect 514587 443816 514789 443817
rect 514587 443616 514588 443816
rect 514788 443616 514789 443816
rect 514587 443615 514789 443616
rect 514587 443416 514789 443417
rect 514587 443216 514588 443416
rect 514788 443216 514789 443416
rect 514587 443215 514789 443216
rect 514587 443016 514789 443017
rect 514587 442816 514588 443016
rect 514788 442816 514789 443016
rect 514587 442815 514789 442816
rect 514587 442616 514789 442617
rect 514587 442416 514588 442616
rect 514788 442416 514789 442616
rect 514587 442415 514789 442416
rect 514587 442216 514789 442217
rect 514587 442016 514588 442216
rect 514788 442016 514789 442216
rect 514587 442015 514789 442016
rect 514587 441816 514789 441817
rect 514587 441616 514588 441816
rect 514788 441616 514789 441816
rect 514587 441615 514789 441616
rect 514587 441416 514789 441417
rect 514587 441216 514588 441416
rect 514788 441216 514789 441416
rect 514587 441215 514789 441216
rect 514587 441016 514789 441017
rect 514587 440816 514588 441016
rect 514788 440816 514789 441016
rect 514587 440815 514789 440816
rect 512233 439887 513207 439888
rect 490464 431892 491260 436676
rect 497004 431892 497126 436676
rect 490464 426000 497126 431892
rect 500384 437540 501424 437596
rect 500384 437440 500418 437540
rect 500518 437440 500642 437540
rect 500742 437440 500866 437540
rect 500966 437440 501090 437540
rect 501190 437440 501314 437540
rect 501414 437440 501424 437540
rect 500384 437316 501424 437440
rect 500384 437216 500418 437316
rect 500518 437216 500642 437316
rect 500742 437216 500866 437316
rect 500966 437216 501090 437316
rect 501190 437216 501314 437316
rect 501414 437216 501424 437316
rect 500384 437092 501424 437216
rect 500384 436992 500418 437092
rect 500518 436992 500642 437092
rect 500742 436992 500866 437092
rect 500966 436992 501090 437092
rect 501190 436992 501314 437092
rect 501414 436992 501424 437092
rect 500384 436868 501424 436992
rect 500384 436768 500418 436868
rect 500518 436768 500642 436868
rect 500742 436768 500866 436868
rect 500966 436768 501090 436868
rect 501190 436768 501314 436868
rect 501414 436768 501424 436868
rect 500384 436644 501424 436768
rect 500384 436544 500418 436644
rect 500518 436544 500642 436644
rect 500742 436544 500866 436644
rect 500966 436544 501090 436644
rect 501190 436544 501314 436644
rect 501414 436544 501424 436644
rect 500384 436420 501424 436544
rect 500384 436320 500418 436420
rect 500518 436320 500642 436420
rect 500742 436320 500866 436420
rect 500966 436320 501090 436420
rect 501190 436320 501314 436420
rect 501414 436320 501424 436420
rect 500384 436196 501424 436320
rect 500384 436096 500418 436196
rect 500518 436096 500642 436196
rect 500742 436096 500866 436196
rect 500966 436096 501090 436196
rect 501190 436096 501314 436196
rect 501414 436096 501424 436196
rect 500384 435972 501424 436096
rect 500384 435872 500418 435972
rect 500518 435872 500642 435972
rect 500742 435872 500866 435972
rect 500966 435872 501090 435972
rect 501190 435872 501314 435972
rect 501414 435872 501424 435972
rect 500384 435748 501424 435872
rect 500384 435648 500418 435748
rect 500518 435648 500642 435748
rect 500742 435648 500866 435748
rect 500966 435648 501090 435748
rect 501190 435648 501314 435748
rect 501414 435648 501424 435748
rect 500384 435524 501424 435648
rect 500384 435424 500418 435524
rect 500518 435424 500642 435524
rect 500742 435424 500866 435524
rect 500966 435424 501090 435524
rect 501190 435424 501314 435524
rect 501414 435424 501424 435524
rect 500384 435300 501424 435424
rect 500384 435200 500418 435300
rect 500518 435200 500642 435300
rect 500742 435200 500866 435300
rect 500966 435200 501090 435300
rect 501190 435200 501314 435300
rect 501414 435200 501424 435300
rect 500384 435076 501424 435200
rect 500384 434976 500418 435076
rect 500518 434976 500642 435076
rect 500742 434976 500866 435076
rect 500966 434976 501090 435076
rect 501190 434976 501314 435076
rect 501414 434976 501424 435076
rect 500384 434852 501424 434976
rect 500384 434752 500418 434852
rect 500518 434752 500642 434852
rect 500742 434752 500866 434852
rect 500966 434752 501090 434852
rect 501190 434752 501314 434852
rect 501414 434752 501424 434852
rect 500384 434628 501424 434752
rect 500384 434528 500418 434628
rect 500518 434528 500642 434628
rect 500742 434528 500866 434628
rect 500966 434528 501090 434628
rect 501190 434528 501314 434628
rect 501414 434528 501424 434628
rect 500384 434404 501424 434528
rect 500384 434304 500418 434404
rect 500518 434304 500642 434404
rect 500742 434304 500866 434404
rect 500966 434304 501090 434404
rect 501190 434304 501314 434404
rect 501414 434304 501424 434404
rect 500384 434180 501424 434304
rect 500384 434080 500418 434180
rect 500518 434080 500642 434180
rect 500742 434080 500866 434180
rect 500966 434080 501090 434180
rect 501190 434080 501314 434180
rect 501414 434080 501424 434180
rect 500384 433956 501424 434080
rect 500384 433856 500418 433956
rect 500518 433856 500642 433956
rect 500742 433856 500866 433956
rect 500966 433856 501090 433956
rect 501190 433856 501314 433956
rect 501414 433856 501424 433956
rect 500384 433732 501424 433856
rect 500384 433632 500418 433732
rect 500518 433632 500642 433732
rect 500742 433632 500866 433732
rect 500966 433632 501090 433732
rect 501190 433632 501314 433732
rect 501414 433632 501424 433732
rect 500384 433508 501424 433632
rect 500384 433408 500418 433508
rect 500518 433408 500642 433508
rect 500742 433408 500866 433508
rect 500966 433408 501090 433508
rect 501190 433408 501314 433508
rect 501414 433408 501424 433508
rect 500384 433284 501424 433408
rect 500384 433184 500418 433284
rect 500518 433184 500642 433284
rect 500742 433184 500866 433284
rect 500966 433184 501090 433284
rect 501190 433184 501314 433284
rect 501414 433184 501424 433284
rect 500384 433060 501424 433184
rect 500384 432960 500418 433060
rect 500518 432960 500642 433060
rect 500742 432960 500866 433060
rect 500966 432960 501090 433060
rect 501190 432960 501314 433060
rect 501414 432960 501424 433060
rect 500384 432836 501424 432960
rect 500384 432736 500418 432836
rect 500518 432736 500642 432836
rect 500742 432736 500866 432836
rect 500966 432736 501090 432836
rect 501190 432736 501314 432836
rect 501414 432736 501424 432836
rect 500384 432612 501424 432736
rect 500384 432512 500418 432612
rect 500518 432512 500642 432612
rect 500742 432512 500866 432612
rect 500966 432512 501090 432612
rect 501190 432512 501314 432612
rect 501414 432512 501424 432612
rect 500384 432388 501424 432512
rect 500384 432288 500418 432388
rect 500518 432288 500642 432388
rect 500742 432288 500866 432388
rect 500966 432288 501090 432388
rect 501190 432288 501314 432388
rect 501414 432288 501424 432388
rect 500384 432164 501424 432288
rect 500384 432064 500418 432164
rect 500518 432064 500642 432164
rect 500742 432064 500866 432164
rect 500966 432064 501090 432164
rect 501190 432064 501314 432164
rect 501414 432064 501424 432164
rect 500384 431940 501424 432064
rect 500384 431840 500418 431940
rect 500518 431840 500642 431940
rect 500742 431840 500866 431940
rect 500966 431840 501090 431940
rect 501190 431840 501314 431940
rect 501414 431840 501424 431940
rect 500384 431716 501424 431840
rect 500384 431616 500418 431716
rect 500518 431616 500642 431716
rect 500742 431616 500866 431716
rect 500966 431616 501090 431716
rect 501190 431616 501314 431716
rect 501414 431616 501424 431716
rect 500384 431492 501424 431616
rect 500384 431392 500418 431492
rect 500518 431392 500642 431492
rect 500742 431392 500866 431492
rect 500966 431392 501090 431492
rect 501190 431392 501314 431492
rect 501414 431392 501424 431492
rect 500384 431268 501424 431392
rect 500384 431168 500418 431268
rect 500518 431168 500642 431268
rect 500742 431168 500866 431268
rect 500966 431168 501090 431268
rect 501190 431168 501314 431268
rect 501414 431168 501424 431268
rect 500384 431044 501424 431168
rect 527604 437540 528644 437596
rect 527604 437440 527638 437540
rect 527738 437440 527862 437540
rect 527962 437440 528086 437540
rect 528186 437440 528310 437540
rect 528410 437440 528534 437540
rect 528634 437440 528644 437540
rect 527604 437316 528644 437440
rect 527604 437216 527638 437316
rect 527738 437216 527862 437316
rect 527962 437216 528086 437316
rect 528186 437216 528310 437316
rect 528410 437216 528534 437316
rect 528634 437216 528644 437316
rect 527604 437092 528644 437216
rect 527604 436992 527638 437092
rect 527738 436992 527862 437092
rect 527962 436992 528086 437092
rect 528186 436992 528310 437092
rect 528410 436992 528534 437092
rect 528634 436992 528644 437092
rect 527604 436868 528644 436992
rect 527604 436768 527638 436868
rect 527738 436768 527862 436868
rect 527962 436768 528086 436868
rect 528186 436768 528310 436868
rect 528410 436768 528534 436868
rect 528634 436768 528644 436868
rect 527604 436644 528644 436768
rect 527604 436544 527638 436644
rect 527738 436544 527862 436644
rect 527962 436544 528086 436644
rect 528186 436544 528310 436644
rect 528410 436544 528534 436644
rect 528634 436544 528644 436644
rect 527604 436420 528644 436544
rect 527604 436320 527638 436420
rect 527738 436320 527862 436420
rect 527962 436320 528086 436420
rect 528186 436320 528310 436420
rect 528410 436320 528534 436420
rect 528634 436320 528644 436420
rect 527604 436196 528644 436320
rect 527604 436096 527638 436196
rect 527738 436096 527862 436196
rect 527962 436096 528086 436196
rect 528186 436096 528310 436196
rect 528410 436096 528534 436196
rect 528634 436096 528644 436196
rect 527604 435972 528644 436096
rect 527604 435872 527638 435972
rect 527738 435872 527862 435972
rect 527962 435872 528086 435972
rect 528186 435872 528310 435972
rect 528410 435872 528534 435972
rect 528634 435872 528644 435972
rect 527604 435748 528644 435872
rect 527604 435648 527638 435748
rect 527738 435648 527862 435748
rect 527962 435648 528086 435748
rect 528186 435648 528310 435748
rect 528410 435648 528534 435748
rect 528634 435648 528644 435748
rect 527604 435524 528644 435648
rect 527604 435424 527638 435524
rect 527738 435424 527862 435524
rect 527962 435424 528086 435524
rect 528186 435424 528310 435524
rect 528410 435424 528534 435524
rect 528634 435424 528644 435524
rect 527604 435300 528644 435424
rect 527604 435200 527638 435300
rect 527738 435200 527862 435300
rect 527962 435200 528086 435300
rect 528186 435200 528310 435300
rect 528410 435200 528534 435300
rect 528634 435200 528644 435300
rect 527604 435076 528644 435200
rect 527604 434976 527638 435076
rect 527738 434976 527862 435076
rect 527962 434976 528086 435076
rect 528186 434976 528310 435076
rect 528410 434976 528534 435076
rect 528634 434976 528644 435076
rect 527604 434852 528644 434976
rect 527604 434752 527638 434852
rect 527738 434752 527862 434852
rect 527962 434752 528086 434852
rect 528186 434752 528310 434852
rect 528410 434752 528534 434852
rect 528634 434752 528644 434852
rect 527604 434628 528644 434752
rect 527604 434528 527638 434628
rect 527738 434528 527862 434628
rect 527962 434528 528086 434628
rect 528186 434528 528310 434628
rect 528410 434528 528534 434628
rect 528634 434528 528644 434628
rect 527604 434404 528644 434528
rect 527604 434304 527638 434404
rect 527738 434304 527862 434404
rect 527962 434304 528086 434404
rect 528186 434304 528310 434404
rect 528410 434304 528534 434404
rect 528634 434304 528644 434404
rect 527604 434180 528644 434304
rect 527604 434080 527638 434180
rect 527738 434080 527862 434180
rect 527962 434080 528086 434180
rect 528186 434080 528310 434180
rect 528410 434080 528534 434180
rect 528634 434080 528644 434180
rect 527604 433956 528644 434080
rect 527604 433856 527638 433956
rect 527738 433856 527862 433956
rect 527962 433856 528086 433956
rect 528186 433856 528310 433956
rect 528410 433856 528534 433956
rect 528634 433856 528644 433956
rect 527604 433732 528644 433856
rect 527604 433632 527638 433732
rect 527738 433632 527862 433732
rect 527962 433632 528086 433732
rect 528186 433632 528310 433732
rect 528410 433632 528534 433732
rect 528634 433632 528644 433732
rect 527604 433508 528644 433632
rect 527604 433408 527638 433508
rect 527738 433408 527862 433508
rect 527962 433408 528086 433508
rect 528186 433408 528310 433508
rect 528410 433408 528534 433508
rect 528634 433408 528644 433508
rect 527604 433284 528644 433408
rect 527604 433184 527638 433284
rect 527738 433184 527862 433284
rect 527962 433184 528086 433284
rect 528186 433184 528310 433284
rect 528410 433184 528534 433284
rect 528634 433184 528644 433284
rect 527604 433060 528644 433184
rect 527604 432960 527638 433060
rect 527738 432960 527862 433060
rect 527962 432960 528086 433060
rect 528186 432960 528310 433060
rect 528410 432960 528534 433060
rect 528634 432960 528644 433060
rect 527604 432836 528644 432960
rect 527604 432736 527638 432836
rect 527738 432736 527862 432836
rect 527962 432736 528086 432836
rect 528186 432736 528310 432836
rect 528410 432736 528534 432836
rect 528634 432736 528644 432836
rect 527604 432612 528644 432736
rect 527604 432512 527638 432612
rect 527738 432512 527862 432612
rect 527962 432512 528086 432612
rect 528186 432512 528310 432612
rect 528410 432512 528534 432612
rect 528634 432512 528644 432612
rect 527604 432388 528644 432512
rect 527604 432288 527638 432388
rect 527738 432288 527862 432388
rect 527962 432288 528086 432388
rect 528186 432288 528310 432388
rect 528410 432288 528534 432388
rect 528634 432288 528644 432388
rect 527604 432164 528644 432288
rect 527604 432064 527638 432164
rect 527738 432064 527862 432164
rect 527962 432064 528086 432164
rect 528186 432064 528310 432164
rect 528410 432064 528534 432164
rect 528634 432064 528644 432164
rect 527604 431940 528644 432064
rect 527604 431840 527638 431940
rect 527738 431840 527862 431940
rect 527962 431840 528086 431940
rect 528186 431840 528310 431940
rect 528410 431840 528534 431940
rect 528634 431840 528644 431940
rect 527604 431716 528644 431840
rect 527604 431616 527638 431716
rect 527738 431616 527862 431716
rect 527962 431616 528086 431716
rect 528186 431616 528310 431716
rect 528410 431616 528534 431716
rect 528634 431616 528644 431716
rect 527604 431492 528644 431616
rect 527604 431392 527638 431492
rect 527738 431392 527862 431492
rect 527962 431392 528086 431492
rect 528186 431392 528310 431492
rect 528410 431392 528534 431492
rect 528634 431392 528644 431492
rect 527604 431268 528644 431392
rect 527604 431168 527638 431268
rect 527738 431168 527862 431268
rect 527962 431168 528086 431268
rect 528186 431168 528310 431268
rect 528410 431168 528534 431268
rect 528634 431168 528644 431268
rect 500384 430944 500418 431044
rect 500518 430944 500642 431044
rect 500742 430944 500866 431044
rect 500966 430944 501090 431044
rect 501190 430944 501314 431044
rect 501414 430944 501424 431044
rect 500384 430940 501424 430944
rect 503864 431026 510526 431156
rect 500413 430939 500523 430940
rect 500637 430939 500747 430940
rect 500861 430939 500971 430940
rect 501085 430939 501195 430940
rect 501309 430939 501419 430940
rect 490464 421216 491138 426000
rect 496882 421216 497126 426000
rect 490464 411200 497126 421216
rect 503864 430926 503920 431026
rect 504020 430926 504144 431026
rect 504244 430926 504368 431026
rect 504468 430926 504592 431026
rect 504692 430926 504816 431026
rect 504916 430926 505040 431026
rect 505140 430926 505264 431026
rect 505364 430926 505488 431026
rect 505588 430926 505712 431026
rect 505812 430926 505936 431026
rect 506036 430926 506160 431026
rect 506260 430926 506384 431026
rect 506484 430926 506608 431026
rect 506708 430926 506832 431026
rect 506932 430926 507056 431026
rect 507156 430926 507280 431026
rect 507380 430926 507504 431026
rect 507604 430926 507728 431026
rect 507828 430926 507952 431026
rect 508052 430926 508176 431026
rect 508276 430926 508400 431026
rect 508500 430926 508624 431026
rect 508724 430926 508848 431026
rect 508948 430926 509072 431026
rect 509172 430926 509296 431026
rect 509396 430926 509520 431026
rect 509620 430926 509744 431026
rect 509844 430926 509968 431026
rect 510068 430926 510192 431026
rect 510292 430926 510416 431026
rect 510516 430926 510526 431026
rect 503864 430802 510526 430926
rect 503864 430702 503920 430802
rect 504020 430702 504144 430802
rect 504244 430702 504368 430802
rect 504468 430702 504592 430802
rect 504692 430702 504816 430802
rect 504916 430702 505040 430802
rect 505140 430702 505264 430802
rect 505364 430702 505488 430802
rect 505588 430702 505712 430802
rect 505812 430702 505936 430802
rect 506036 430702 506160 430802
rect 506260 430702 506384 430802
rect 506484 430702 506608 430802
rect 506708 430702 506832 430802
rect 506932 430702 507056 430802
rect 507156 430702 507280 430802
rect 507380 430702 507504 430802
rect 507604 430702 507728 430802
rect 507828 430702 507952 430802
rect 508052 430702 508176 430802
rect 508276 430702 508400 430802
rect 508500 430702 508624 430802
rect 508724 430702 508848 430802
rect 508948 430702 509072 430802
rect 509172 430702 509296 430802
rect 509396 430702 509520 430802
rect 509620 430702 509744 430802
rect 509844 430702 509968 430802
rect 510068 430702 510192 430802
rect 510292 430702 510416 430802
rect 510516 430702 510526 430802
rect 503864 430578 510526 430702
rect 503864 430478 503920 430578
rect 504020 430478 504144 430578
rect 504244 430478 504368 430578
rect 504468 430478 504592 430578
rect 504692 430478 504816 430578
rect 504916 430478 505040 430578
rect 505140 430478 505264 430578
rect 505364 430478 505488 430578
rect 505588 430478 505712 430578
rect 505812 430478 505936 430578
rect 506036 430478 506160 430578
rect 506260 430478 506384 430578
rect 506484 430478 506608 430578
rect 506708 430478 506832 430578
rect 506932 430478 507056 430578
rect 507156 430478 507280 430578
rect 507380 430478 507504 430578
rect 507604 430478 507728 430578
rect 507828 430478 507952 430578
rect 508052 430478 508176 430578
rect 508276 430478 508400 430578
rect 508500 430478 508624 430578
rect 508724 430478 508848 430578
rect 508948 430478 509072 430578
rect 509172 430478 509296 430578
rect 509396 430478 509520 430578
rect 509620 430478 509744 430578
rect 509844 430478 509968 430578
rect 510068 430478 510192 430578
rect 510292 430478 510416 430578
rect 510516 430478 510526 430578
rect 503864 430354 510526 430478
rect 503864 430254 503920 430354
rect 504020 430254 504144 430354
rect 504244 430254 504368 430354
rect 504468 430254 504592 430354
rect 504692 430254 504816 430354
rect 504916 430254 505040 430354
rect 505140 430254 505264 430354
rect 505364 430254 505488 430354
rect 505588 430254 505712 430354
rect 505812 430254 505936 430354
rect 506036 430254 506160 430354
rect 506260 430254 506384 430354
rect 506484 430254 506608 430354
rect 506708 430254 506832 430354
rect 506932 430254 507056 430354
rect 507156 430254 507280 430354
rect 507380 430254 507504 430354
rect 507604 430254 507728 430354
rect 507828 430254 507952 430354
rect 508052 430254 508176 430354
rect 508276 430254 508400 430354
rect 508500 430254 508624 430354
rect 508724 430254 508848 430354
rect 508948 430254 509072 430354
rect 509172 430254 509296 430354
rect 509396 430254 509520 430354
rect 509620 430254 509744 430354
rect 509844 430254 509968 430354
rect 510068 430254 510192 430354
rect 510292 430254 510416 430354
rect 510516 430254 510526 430354
rect 503864 430130 510526 430254
rect 503864 430030 503920 430130
rect 504020 430030 504144 430130
rect 504244 430030 504368 430130
rect 504468 430030 504592 430130
rect 504692 430030 504816 430130
rect 504916 430030 505040 430130
rect 505140 430030 505264 430130
rect 505364 430030 505488 430130
rect 505588 430030 505712 430130
rect 505812 430030 505936 430130
rect 506036 430030 506160 430130
rect 506260 430030 506384 430130
rect 506484 430030 506608 430130
rect 506708 430030 506832 430130
rect 506932 430030 507056 430130
rect 507156 430030 507280 430130
rect 507380 430030 507504 430130
rect 507604 430030 507728 430130
rect 507828 430030 507952 430130
rect 508052 430030 508176 430130
rect 508276 430030 508400 430130
rect 508500 430030 508624 430130
rect 508724 430030 508848 430130
rect 508948 430030 509072 430130
rect 509172 430030 509296 430130
rect 509396 430030 509520 430130
rect 509620 430030 509744 430130
rect 509844 430030 509968 430130
rect 510068 430030 510192 430130
rect 510292 430030 510416 430130
rect 510516 430030 510526 430130
rect 503864 426000 510526 430030
rect 503864 421216 504338 426000
rect 510082 421216 510526 426000
rect 503864 420526 510526 421216
rect 517264 431031 523920 431162
rect 527604 431044 528644 431168
rect 517264 431026 523921 431031
rect 517264 430926 517320 431026
rect 517420 430926 517544 431026
rect 517644 430926 517768 431026
rect 517868 430926 517992 431026
rect 518092 430926 518216 431026
rect 518316 430926 518440 431026
rect 518540 430926 518664 431026
rect 518764 430926 518888 431026
rect 518988 430926 519112 431026
rect 519212 430926 519336 431026
rect 519436 430926 519560 431026
rect 519660 430926 519784 431026
rect 519884 430926 520008 431026
rect 520108 430926 520232 431026
rect 520332 430926 520456 431026
rect 520556 430926 520680 431026
rect 520780 430926 520904 431026
rect 521004 430926 521128 431026
rect 521228 430926 521352 431026
rect 521452 430926 521576 431026
rect 521676 430926 521800 431026
rect 521900 430926 522024 431026
rect 522124 430926 522248 431026
rect 522348 430926 522472 431026
rect 522572 430926 522696 431026
rect 522796 430926 522920 431026
rect 523020 430926 523144 431026
rect 523244 430926 523368 431026
rect 523468 430926 523592 431026
rect 523692 430926 523816 431026
rect 523916 430926 523921 431026
rect 527604 430944 527638 431044
rect 527738 430944 527862 431044
rect 527962 430944 528086 431044
rect 528186 430944 528310 431044
rect 528410 430944 528534 431044
rect 528634 430944 528644 431044
rect 527604 430940 528644 430944
rect 530664 436676 537320 457452
rect 562380 455480 567480 455520
rect 562380 455440 562624 455480
rect 562860 455440 563096 455480
rect 563332 455440 563568 455480
rect 563804 455440 564040 455480
rect 564276 455440 564512 455480
rect 564748 455440 564984 455480
rect 565220 455440 565456 455480
rect 565692 455440 565928 455480
rect 566164 455440 566400 455480
rect 566636 455440 566872 455480
rect 567108 455440 567480 455480
rect 562380 455360 562480 455440
rect 562560 455360 562624 455440
rect 562880 455360 562960 455440
rect 563040 455360 563096 455440
rect 563360 455360 563440 455440
rect 563520 455360 563568 455440
rect 563840 455360 563920 455440
rect 564000 455360 564040 455440
rect 564320 455360 564400 455440
rect 564480 455360 564512 455440
rect 564800 455360 564880 455440
rect 564960 455360 564984 455440
rect 565280 455360 565360 455440
rect 565440 455360 565456 455440
rect 565760 455360 565840 455440
rect 565920 455360 565928 455440
rect 566240 455360 566320 455440
rect 566636 455360 566640 455440
rect 566720 455360 566800 455440
rect 567108 455360 567120 455440
rect 567200 455360 567280 455440
rect 567360 455360 567480 455440
rect 562380 455280 562624 455360
rect 562860 455280 563096 455360
rect 563332 455280 563568 455360
rect 563804 455280 564040 455360
rect 564276 455280 564512 455360
rect 564748 455280 564984 455360
rect 565220 455280 565456 455360
rect 565692 455280 565928 455360
rect 566164 455280 566400 455360
rect 566636 455280 566872 455360
rect 567108 455280 567480 455360
rect 562380 455200 562480 455280
rect 562560 455244 562624 455280
rect 562560 455200 562640 455244
rect 562720 455200 562800 455244
rect 562880 455200 562960 455280
rect 563040 455244 563096 455280
rect 563040 455200 563120 455244
rect 563200 455200 563280 455244
rect 563360 455200 563440 455280
rect 563520 455244 563568 455280
rect 563520 455200 563600 455244
rect 563680 455200 563760 455244
rect 563840 455200 563920 455280
rect 564000 455244 564040 455280
rect 564000 455200 564080 455244
rect 564160 455200 564240 455244
rect 564320 455200 564400 455280
rect 564480 455244 564512 455280
rect 564480 455200 564560 455244
rect 564640 455200 564720 455244
rect 564800 455200 564880 455280
rect 564960 455244 564984 455280
rect 564960 455200 565040 455244
rect 565120 455200 565200 455244
rect 565280 455200 565360 455280
rect 565440 455244 565456 455280
rect 565440 455200 565520 455244
rect 565600 455200 565680 455244
rect 565760 455200 565840 455280
rect 565920 455244 565928 455280
rect 565920 455200 566000 455244
rect 566080 455200 566160 455244
rect 566240 455200 566320 455280
rect 566636 455244 566640 455280
rect 566400 455200 566480 455244
rect 566560 455200 566640 455244
rect 566720 455200 566800 455280
rect 567108 455244 567120 455280
rect 566880 455200 566960 455244
rect 567040 455200 567120 455244
rect 567200 455200 567280 455280
rect 567360 455200 567480 455280
rect 562380 455160 567480 455200
rect 572540 455480 577640 455520
rect 572540 455440 572784 455480
rect 573020 455440 573256 455480
rect 573492 455440 573728 455480
rect 573964 455440 574200 455480
rect 574436 455440 574672 455480
rect 574908 455440 575144 455480
rect 575380 455440 575616 455480
rect 575852 455440 576088 455480
rect 576324 455440 576560 455480
rect 576796 455440 577032 455480
rect 577268 455440 577640 455480
rect 572540 455360 572640 455440
rect 572720 455360 572784 455440
rect 573040 455360 573120 455440
rect 573200 455360 573256 455440
rect 573520 455360 573600 455440
rect 573680 455360 573728 455440
rect 574000 455360 574080 455440
rect 574160 455360 574200 455440
rect 574480 455360 574560 455440
rect 574640 455360 574672 455440
rect 574960 455360 575040 455440
rect 575120 455360 575144 455440
rect 575440 455360 575520 455440
rect 575600 455360 575616 455440
rect 575920 455360 576000 455440
rect 576080 455360 576088 455440
rect 576400 455360 576480 455440
rect 576796 455360 576800 455440
rect 576880 455360 576960 455440
rect 577268 455360 577280 455440
rect 577360 455360 577440 455440
rect 577520 455360 577640 455440
rect 572540 455280 572784 455360
rect 573020 455280 573256 455360
rect 573492 455280 573728 455360
rect 573964 455280 574200 455360
rect 574436 455280 574672 455360
rect 574908 455280 575144 455360
rect 575380 455280 575616 455360
rect 575852 455280 576088 455360
rect 576324 455280 576560 455360
rect 576796 455280 577032 455360
rect 577268 455280 577640 455360
rect 572540 455200 572640 455280
rect 572720 455244 572784 455280
rect 572720 455200 572800 455244
rect 572880 455200 572960 455244
rect 573040 455200 573120 455280
rect 573200 455244 573256 455280
rect 573200 455200 573280 455244
rect 573360 455200 573440 455244
rect 573520 455200 573600 455280
rect 573680 455244 573728 455280
rect 573680 455200 573760 455244
rect 573840 455200 573920 455244
rect 574000 455200 574080 455280
rect 574160 455244 574200 455280
rect 574160 455200 574240 455244
rect 574320 455200 574400 455244
rect 574480 455200 574560 455280
rect 574640 455244 574672 455280
rect 574640 455200 574720 455244
rect 574800 455200 574880 455244
rect 574960 455200 575040 455280
rect 575120 455244 575144 455280
rect 575120 455200 575200 455244
rect 575280 455200 575360 455244
rect 575440 455200 575520 455280
rect 575600 455244 575616 455280
rect 575600 455200 575680 455244
rect 575760 455200 575840 455244
rect 575920 455200 576000 455280
rect 576080 455244 576088 455280
rect 576080 455200 576160 455244
rect 576240 455200 576320 455244
rect 576400 455200 576480 455280
rect 576796 455244 576800 455280
rect 576560 455200 576640 455244
rect 576720 455200 576800 455244
rect 576880 455200 576960 455280
rect 577268 455244 577280 455280
rect 577040 455200 577120 455244
rect 577200 455200 577280 455244
rect 577360 455200 577440 455280
rect 577520 455200 577640 455280
rect 572540 455160 577640 455200
rect 530664 431892 531080 436676
rect 536824 431892 537320 436676
rect 527633 430939 527743 430940
rect 527857 430939 527967 430940
rect 528081 430939 528191 430940
rect 528305 430939 528415 430940
rect 528529 430939 528639 430940
rect 517264 430921 523921 430926
rect 517264 430807 523920 430921
rect 517264 430802 523921 430807
rect 517264 430702 517320 430802
rect 517420 430702 517544 430802
rect 517644 430702 517768 430802
rect 517868 430702 517992 430802
rect 518092 430702 518216 430802
rect 518316 430702 518440 430802
rect 518540 430702 518664 430802
rect 518764 430702 518888 430802
rect 518988 430702 519112 430802
rect 519212 430702 519336 430802
rect 519436 430702 519560 430802
rect 519660 430702 519784 430802
rect 519884 430702 520008 430802
rect 520108 430702 520232 430802
rect 520332 430702 520456 430802
rect 520556 430702 520680 430802
rect 520780 430702 520904 430802
rect 521004 430702 521128 430802
rect 521228 430702 521352 430802
rect 521452 430702 521576 430802
rect 521676 430702 521800 430802
rect 521900 430702 522024 430802
rect 522124 430702 522248 430802
rect 522348 430702 522472 430802
rect 522572 430702 522696 430802
rect 522796 430702 522920 430802
rect 523020 430702 523144 430802
rect 523244 430702 523368 430802
rect 523468 430702 523592 430802
rect 523692 430702 523816 430802
rect 523916 430702 523921 430802
rect 517264 430697 523921 430702
rect 517264 430583 523920 430697
rect 517264 430578 523921 430583
rect 517264 430478 517320 430578
rect 517420 430478 517544 430578
rect 517644 430478 517768 430578
rect 517868 430478 517992 430578
rect 518092 430478 518216 430578
rect 518316 430478 518440 430578
rect 518540 430478 518664 430578
rect 518764 430478 518888 430578
rect 518988 430478 519112 430578
rect 519212 430478 519336 430578
rect 519436 430478 519560 430578
rect 519660 430478 519784 430578
rect 519884 430478 520008 430578
rect 520108 430478 520232 430578
rect 520332 430478 520456 430578
rect 520556 430478 520680 430578
rect 520780 430478 520904 430578
rect 521004 430478 521128 430578
rect 521228 430478 521352 430578
rect 521452 430478 521576 430578
rect 521676 430478 521800 430578
rect 521900 430478 522024 430578
rect 522124 430478 522248 430578
rect 522348 430478 522472 430578
rect 522572 430478 522696 430578
rect 522796 430478 522920 430578
rect 523020 430478 523144 430578
rect 523244 430478 523368 430578
rect 523468 430478 523592 430578
rect 523692 430478 523816 430578
rect 523916 430478 523921 430578
rect 517264 430473 523921 430478
rect 517264 430359 523920 430473
rect 517264 430354 523921 430359
rect 517264 430254 517320 430354
rect 517420 430254 517544 430354
rect 517644 430254 517768 430354
rect 517868 430254 517992 430354
rect 518092 430254 518216 430354
rect 518316 430254 518440 430354
rect 518540 430254 518664 430354
rect 518764 430254 518888 430354
rect 518988 430254 519112 430354
rect 519212 430254 519336 430354
rect 519436 430254 519560 430354
rect 519660 430254 519784 430354
rect 519884 430254 520008 430354
rect 520108 430254 520232 430354
rect 520332 430254 520456 430354
rect 520556 430254 520680 430354
rect 520780 430254 520904 430354
rect 521004 430254 521128 430354
rect 521228 430254 521352 430354
rect 521452 430254 521576 430354
rect 521676 430254 521800 430354
rect 521900 430254 522024 430354
rect 522124 430254 522248 430354
rect 522348 430254 522472 430354
rect 522572 430254 522696 430354
rect 522796 430254 522920 430354
rect 523020 430254 523144 430354
rect 523244 430254 523368 430354
rect 523468 430254 523592 430354
rect 523692 430254 523816 430354
rect 523916 430254 523921 430354
rect 517264 430249 523921 430254
rect 517264 430135 523920 430249
rect 517264 430130 523921 430135
rect 517264 430030 517320 430130
rect 517420 430030 517544 430130
rect 517644 430030 517768 430130
rect 517868 430030 517992 430130
rect 518092 430030 518216 430130
rect 518316 430030 518440 430130
rect 518540 430030 518664 430130
rect 518764 430030 518888 430130
rect 518988 430030 519112 430130
rect 519212 430030 519336 430130
rect 519436 430030 519560 430130
rect 519660 430030 519784 430130
rect 519884 430030 520008 430130
rect 520108 430030 520232 430130
rect 520332 430030 520456 430130
rect 520556 430030 520680 430130
rect 520780 430030 520904 430130
rect 521004 430030 521128 430130
rect 521228 430030 521352 430130
rect 521452 430030 521576 430130
rect 521676 430030 521800 430130
rect 521900 430030 522024 430130
rect 522124 430030 522248 430130
rect 522348 430030 522472 430130
rect 522572 430030 522696 430130
rect 522796 430030 522920 430130
rect 523020 430030 523144 430130
rect 523244 430030 523368 430130
rect 523468 430030 523592 430130
rect 523692 430030 523816 430130
rect 523916 430030 523921 430130
rect 517264 430025 523921 430030
rect 517264 426000 523920 430025
rect 517264 421216 517738 426000
rect 523482 421216 523920 426000
rect 517264 420526 523920 421216
rect 530664 429736 537320 431892
rect 530664 426000 537326 429736
rect 530664 421216 531138 426000
rect 536882 425278 537326 426000
rect 572536 426688 577492 426924
rect 536882 421216 537320 425278
rect 530664 415278 537320 421216
rect 572536 420316 572772 426688
rect 573008 420316 573244 426688
rect 573480 420316 573716 426688
rect 573952 420316 574188 426688
rect 574424 420316 574660 426688
rect 574896 420316 575132 426688
rect 575368 420316 575604 426688
rect 575840 420316 576076 426688
rect 576312 420316 576548 426688
rect 576784 420316 577020 426688
rect 577256 420316 577492 426688
rect 477060 377836 483800 378072
rect 477060 377600 477192 377836
rect 477428 377600 477664 377836
rect 477900 377600 478136 377836
rect 478372 377600 478608 377836
rect 478844 377600 479080 377836
rect 479316 377600 479552 377836
rect 479788 377600 480024 377836
rect 480260 377600 480496 377836
rect 480732 377600 480968 377836
rect 481204 377600 481440 377836
rect 481676 377600 481912 377836
rect 482148 377600 482384 377836
rect 482620 377600 482856 377836
rect 483092 377600 483328 377836
rect 483564 377600 483800 377836
rect 477060 377364 483800 377600
rect 477060 377128 477192 377364
rect 477428 377128 477664 377364
rect 477900 377128 478136 377364
rect 478372 377128 478608 377364
rect 478844 377128 479080 377364
rect 479316 377128 479552 377364
rect 479788 377128 480024 377364
rect 480260 377128 480496 377364
rect 480732 377128 480968 377364
rect 481204 377128 481440 377364
rect 481676 377128 481912 377364
rect 482148 377128 482384 377364
rect 482620 377128 482856 377364
rect 483092 377128 483328 377364
rect 483564 377128 483800 377364
rect 477060 376892 483800 377128
rect 477060 376656 477192 376892
rect 477428 376656 477664 376892
rect 477900 376656 478136 376892
rect 478372 376656 478608 376892
rect 478844 376656 479080 376892
rect 479316 376656 479552 376892
rect 479788 376656 480024 376892
rect 480260 376656 480496 376892
rect 480732 376656 480968 376892
rect 481204 376656 481440 376892
rect 481676 376656 481912 376892
rect 482148 376656 482384 376892
rect 482620 376656 482856 376892
rect 483092 376656 483328 376892
rect 483564 376656 483800 376892
rect 477060 376420 483800 376656
rect 477060 376184 477192 376420
rect 477428 376184 477664 376420
rect 477900 376184 478136 376420
rect 478372 376184 478608 376420
rect 478844 376184 479080 376420
rect 479316 376184 479552 376420
rect 479788 376184 480024 376420
rect 480260 376184 480496 376420
rect 480732 376184 480968 376420
rect 481204 376184 481440 376420
rect 481676 376184 481912 376420
rect 482148 376184 482384 376420
rect 482620 376184 482856 376420
rect 483092 376184 483328 376420
rect 483564 376184 483800 376420
rect 477060 375948 483800 376184
rect 477060 375712 477192 375948
rect 477428 375712 477664 375948
rect 477900 375712 478136 375948
rect 478372 375712 478608 375948
rect 478844 375712 479080 375948
rect 479316 375712 479552 375948
rect 479788 375712 480024 375948
rect 480260 375712 480496 375948
rect 480732 375712 480968 375948
rect 481204 375712 481440 375948
rect 481676 375712 481912 375948
rect 482148 375712 482384 375948
rect 482620 375712 482856 375948
rect 483092 375712 483328 375948
rect 483564 375712 483800 375948
rect 477060 375476 483800 375712
rect 477060 375240 477192 375476
rect 477428 375240 477664 375476
rect 477900 375240 478136 375476
rect 478372 375240 478608 375476
rect 478844 375240 479080 375476
rect 479316 375240 479552 375476
rect 479788 375240 480024 375476
rect 480260 375240 480496 375476
rect 480732 375240 480968 375476
rect 481204 375240 481440 375476
rect 481676 375240 481912 375476
rect 482148 375240 482384 375476
rect 482620 375240 482856 375476
rect 483092 375240 483328 375476
rect 483564 375240 483800 375476
rect 477060 375004 483800 375240
rect 477060 374768 477192 375004
rect 477428 374768 477664 375004
rect 477900 374768 478136 375004
rect 478372 374768 478608 375004
rect 478844 374768 479080 375004
rect 479316 374768 479552 375004
rect 479788 374768 480024 375004
rect 480260 374768 480496 375004
rect 480732 374768 480968 375004
rect 481204 374768 481440 375004
rect 481676 374768 481912 375004
rect 482148 374768 482384 375004
rect 482620 374768 482856 375004
rect 483092 374768 483328 375004
rect 483564 374768 483800 375004
rect 477060 374532 483800 374768
rect 477060 374296 477192 374532
rect 477428 374296 477664 374532
rect 477900 374296 478136 374532
rect 478372 374296 478608 374532
rect 478844 374296 479080 374532
rect 479316 374296 479552 374532
rect 479788 374296 480024 374532
rect 480260 374296 480496 374532
rect 480732 374296 480968 374532
rect 481204 374296 481440 374532
rect 481676 374296 481912 374532
rect 482148 374296 482384 374532
rect 482620 374296 482856 374532
rect 483092 374296 483328 374532
rect 483564 374296 483800 374532
rect 477060 374060 483800 374296
rect 477060 373824 477192 374060
rect 477428 373824 477664 374060
rect 477900 373824 478136 374060
rect 478372 373824 478608 374060
rect 478844 373824 479080 374060
rect 479316 373824 479552 374060
rect 479788 373824 480024 374060
rect 480260 373824 480496 374060
rect 480732 373824 480968 374060
rect 481204 373824 481440 374060
rect 481676 373824 481912 374060
rect 482148 373824 482384 374060
rect 482620 373824 482856 374060
rect 483092 373824 483328 374060
rect 483564 373824 483800 374060
rect 477060 373588 483800 373824
rect 477060 373352 477192 373588
rect 477428 373352 477664 373588
rect 477900 373352 478136 373588
rect 478372 373352 478608 373588
rect 478844 373352 479080 373588
rect 479316 373352 479552 373588
rect 479788 373352 480024 373588
rect 480260 373352 480496 373588
rect 480732 373352 480968 373588
rect 481204 373352 481440 373588
rect 481676 373352 481912 373588
rect 482148 373352 482384 373588
rect 482620 373352 482856 373588
rect 483092 373352 483328 373588
rect 483564 373352 483800 373588
rect 477060 373116 483800 373352
rect 477060 372880 477192 373116
rect 477428 372880 477664 373116
rect 477900 372880 478136 373116
rect 478372 372880 478608 373116
rect 478844 372880 479080 373116
rect 479316 372880 479552 373116
rect 479788 372880 480024 373116
rect 480260 372880 480496 373116
rect 480732 372880 480968 373116
rect 481204 372880 481440 373116
rect 481676 372880 481912 373116
rect 482148 372880 482384 373116
rect 482620 372880 482856 373116
rect 483092 372880 483328 373116
rect 483564 372880 483800 373116
rect 477060 372644 483800 372880
rect 477060 372408 477192 372644
rect 477428 372408 477664 372644
rect 477900 372408 478136 372644
rect 478372 372408 478608 372644
rect 478844 372408 479080 372644
rect 479316 372408 479552 372644
rect 479788 372408 480024 372644
rect 480260 372408 480496 372644
rect 480732 372408 480968 372644
rect 481204 372408 481440 372644
rect 481676 372408 481912 372644
rect 482148 372408 482384 372644
rect 482620 372408 482856 372644
rect 483092 372408 483328 372644
rect 483564 372408 483800 372644
rect 477060 372172 483800 372408
rect 477060 371936 477192 372172
rect 477428 371936 477664 372172
rect 477900 371936 478136 372172
rect 478372 371936 478608 372172
rect 478844 371936 479080 372172
rect 479316 371936 479552 372172
rect 479788 371936 480024 372172
rect 480260 371936 480496 372172
rect 480732 371936 480968 372172
rect 481204 371936 481440 372172
rect 481676 371936 481912 372172
rect 482148 371936 482384 372172
rect 482620 371936 482856 372172
rect 483092 371936 483328 372172
rect 483564 371936 483800 372172
rect 477060 371700 483800 371936
rect 477060 371464 477192 371700
rect 477428 371464 477664 371700
rect 477900 371464 478136 371700
rect 478372 371464 478608 371700
rect 478844 371464 479080 371700
rect 479316 371464 479552 371700
rect 479788 371464 480024 371700
rect 480260 371464 480496 371700
rect 480732 371464 480968 371700
rect 481204 371464 481440 371700
rect 481676 371464 481912 371700
rect 482148 371464 482384 371700
rect 482620 371464 482856 371700
rect 483092 371464 483328 371700
rect 483564 371464 483800 371700
rect 562388 377600 567816 378072
rect 477060 371200 483726 371464
rect 562388 371228 562624 377600
rect 562860 371228 563096 377600
rect 563332 371228 563568 377600
rect 563804 371228 564040 377600
rect 564276 371228 564512 377600
rect 564748 371228 564984 377600
rect 565220 371228 565456 377600
rect 565692 371228 565928 377600
rect 566164 371228 566400 377600
rect 566636 371228 566872 377600
rect 567108 371228 567816 377600
rect 562388 370992 567816 371228
<< via4 >>
rect 572772 696908 573008 697144
rect 573244 696908 573480 697144
rect 573716 696908 573952 697144
rect 574188 696908 574424 697144
rect 574660 696908 574896 697144
rect 575132 696908 575368 697144
rect 575604 696908 575840 697144
rect 576076 696908 576312 697144
rect 576548 696908 576784 697144
rect 577020 696908 577256 697144
rect 572772 696436 573008 696672
rect 573244 696436 573480 696672
rect 573716 696436 573952 696672
rect 574188 696436 574424 696672
rect 574660 696436 574896 696672
rect 575132 696436 575368 696672
rect 575604 696436 575840 696672
rect 576076 696436 576312 696672
rect 576548 696436 576784 696672
rect 577020 696436 577256 696672
rect 572772 695964 573008 696200
rect 573244 695964 573480 696200
rect 573716 695964 573952 696200
rect 574188 695964 574424 696200
rect 574660 695964 574896 696200
rect 575132 695964 575368 696200
rect 575604 695964 575840 696200
rect 576076 695964 576312 696200
rect 576548 695964 576784 696200
rect 577020 695964 577256 696200
rect 572772 695492 573008 695728
rect 573244 695492 573480 695728
rect 573716 695492 573952 695728
rect 574188 695492 574424 695728
rect 574660 695492 574896 695728
rect 575132 695492 575368 695728
rect 575604 695492 575840 695728
rect 576076 695492 576312 695728
rect 576548 695492 576784 695728
rect 577020 695492 577256 695728
rect 572772 695020 573008 695256
rect 573244 695020 573480 695256
rect 573716 695020 573952 695256
rect 574188 695020 574424 695256
rect 574660 695020 574896 695256
rect 575132 695020 575368 695256
rect 575604 695020 575840 695256
rect 576076 695020 576312 695256
rect 576548 695020 576784 695256
rect 577020 695020 577256 695256
rect 572772 694548 573008 694784
rect 573244 694548 573480 694784
rect 573716 694548 573952 694784
rect 574188 694548 574424 694784
rect 574660 694548 574896 694784
rect 575132 694548 575368 694784
rect 575604 694548 575840 694784
rect 576076 694548 576312 694784
rect 576548 694548 576784 694784
rect 577020 694548 577256 694784
rect 572772 694076 573008 694312
rect 573244 694076 573480 694312
rect 573716 694076 573952 694312
rect 574188 694076 574424 694312
rect 574660 694076 574896 694312
rect 575132 694076 575368 694312
rect 575604 694076 575840 694312
rect 576076 694076 576312 694312
rect 576548 694076 576784 694312
rect 577020 694076 577256 694312
rect 572772 693604 573008 693840
rect 573244 693604 573480 693840
rect 573716 693604 573952 693840
rect 574188 693604 574424 693840
rect 574660 693604 574896 693840
rect 575132 693604 575368 693840
rect 575604 693604 575840 693840
rect 576076 693604 576312 693840
rect 576548 693604 576784 693840
rect 577020 693604 577256 693840
rect 572772 693132 573008 693368
rect 573244 693132 573480 693368
rect 573716 693132 573952 693368
rect 574188 693132 574424 693368
rect 574660 693132 574896 693368
rect 575132 693132 575368 693368
rect 575604 693132 575840 693368
rect 576076 693132 576312 693368
rect 576548 693132 576784 693368
rect 577020 693132 577256 693368
rect 572772 692660 573008 692896
rect 573244 692660 573480 692896
rect 573716 692660 573952 692896
rect 574188 692660 574424 692896
rect 574660 692660 574896 692896
rect 575132 692660 575368 692896
rect 575604 692660 575840 692896
rect 576076 692660 576312 692896
rect 576548 692660 576784 692896
rect 577020 692660 577256 692896
rect 562480 644524 567400 644584
rect 562480 639844 562600 644524
rect 562600 639844 567400 644524
rect 562480 639784 567400 639844
rect 562480 634524 567400 634584
rect 562480 629844 562600 634524
rect 562600 629844 567400 634524
rect 562480 629784 567400 629844
rect 562624 522268 562860 522504
rect 562624 521796 562860 522032
rect 562624 521324 562860 521560
rect 562624 520852 562860 521088
rect 562624 520380 562860 520616
rect 562624 519908 562860 520144
rect 562624 519436 562860 519672
rect 562624 518964 562860 519200
rect 562624 518492 562860 518728
rect 562624 518020 562860 518256
rect 562624 517548 562860 517784
rect 562624 517076 562860 517312
rect 562624 516604 562860 516840
rect 563096 522268 563332 522504
rect 563096 521796 563332 522032
rect 563096 521324 563332 521560
rect 563096 520852 563332 521088
rect 563096 520380 563332 520616
rect 563096 519908 563332 520144
rect 563096 519436 563332 519672
rect 563096 518964 563332 519200
rect 563096 518492 563332 518728
rect 563096 518020 563332 518256
rect 563096 517548 563332 517784
rect 563096 517076 563332 517312
rect 563096 516604 563332 516840
rect 563568 522268 563804 522504
rect 563568 521796 563804 522032
rect 563568 521324 563804 521560
rect 563568 520852 563804 521088
rect 563568 520380 563804 520616
rect 563568 519908 563804 520144
rect 563568 519436 563804 519672
rect 563568 518964 563804 519200
rect 563568 518492 563804 518728
rect 563568 518020 563804 518256
rect 563568 517548 563804 517784
rect 563568 517076 563804 517312
rect 563568 516604 563804 516840
rect 564040 522268 564276 522504
rect 564040 521796 564276 522032
rect 564040 521324 564276 521560
rect 564040 520852 564276 521088
rect 564040 520380 564276 520616
rect 564040 519908 564276 520144
rect 564040 519436 564276 519672
rect 564040 518964 564276 519200
rect 564040 518492 564276 518728
rect 564040 518020 564276 518256
rect 564040 517548 564276 517784
rect 564040 517076 564276 517312
rect 564040 516604 564276 516840
rect 564512 522268 564748 522504
rect 564512 521796 564748 522032
rect 564512 521324 564748 521560
rect 564512 520852 564748 521088
rect 564512 520380 564748 520616
rect 564512 519908 564748 520144
rect 564512 519436 564748 519672
rect 564512 518964 564748 519200
rect 564512 518492 564748 518728
rect 564512 518020 564748 518256
rect 564512 517548 564748 517784
rect 564512 517076 564748 517312
rect 564512 516604 564748 516840
rect 564984 522268 565220 522504
rect 564984 521796 565220 522032
rect 564984 521324 565220 521560
rect 564984 520852 565220 521088
rect 564984 520380 565220 520616
rect 564984 519908 565220 520144
rect 564984 519436 565220 519672
rect 564984 518964 565220 519200
rect 564984 518492 565220 518728
rect 564984 518020 565220 518256
rect 564984 517548 565220 517784
rect 564984 517076 565220 517312
rect 564984 516604 565220 516840
rect 565456 522268 565692 522504
rect 565456 521796 565692 522032
rect 565456 521324 565692 521560
rect 565456 520852 565692 521088
rect 565456 520380 565692 520616
rect 565456 519908 565692 520144
rect 565456 519436 565692 519672
rect 565456 518964 565692 519200
rect 565456 518492 565692 518728
rect 565456 518020 565692 518256
rect 565456 517548 565692 517784
rect 565456 517076 565692 517312
rect 565456 516604 565692 516840
rect 565928 522268 566164 522504
rect 565928 521796 566164 522032
rect 565928 521324 566164 521560
rect 565928 520852 566164 521088
rect 565928 520380 566164 520616
rect 565928 519908 566164 520144
rect 565928 519436 566164 519672
rect 565928 518964 566164 519200
rect 565928 518492 566164 518728
rect 565928 518020 566164 518256
rect 565928 517548 566164 517784
rect 565928 517076 566164 517312
rect 565928 516604 566164 516840
rect 566400 522268 566636 522504
rect 566400 521796 566636 522032
rect 566400 521324 566636 521560
rect 566400 520852 566636 521088
rect 566400 520380 566636 520616
rect 566400 519908 566636 520144
rect 566400 519436 566636 519672
rect 566400 518964 566636 519200
rect 566400 518492 566636 518728
rect 566400 518020 566636 518256
rect 566400 517548 566636 517784
rect 566400 517076 566636 517312
rect 566400 516604 566636 516840
rect 566872 522268 567108 522504
rect 566872 521796 567108 522032
rect 566872 521324 567108 521560
rect 566872 520852 567108 521088
rect 566872 520380 567108 520616
rect 566872 519908 567108 520144
rect 566872 519436 567108 519672
rect 566872 518964 567108 519200
rect 566872 518492 567108 518728
rect 566872 518020 567108 518256
rect 566872 517548 567108 517784
rect 566872 517076 567108 517312
rect 566872 516604 567108 516840
rect 562624 495742 562860 495782
rect 563096 495742 563332 495782
rect 563568 495742 563804 495782
rect 564040 495742 564276 495782
rect 564512 495742 564748 495782
rect 564984 495742 565220 495782
rect 565456 495742 565692 495782
rect 565928 495742 566164 495782
rect 566400 495742 566636 495782
rect 566872 495742 567108 495782
rect 562624 495662 562640 495742
rect 562640 495662 562720 495742
rect 562720 495662 562800 495742
rect 562800 495662 562860 495742
rect 563096 495662 563120 495742
rect 563120 495662 563200 495742
rect 563200 495662 563280 495742
rect 563280 495662 563332 495742
rect 563568 495662 563600 495742
rect 563600 495662 563680 495742
rect 563680 495662 563760 495742
rect 563760 495662 563804 495742
rect 564040 495662 564080 495742
rect 564080 495662 564160 495742
rect 564160 495662 564240 495742
rect 564240 495662 564276 495742
rect 564512 495662 564560 495742
rect 564560 495662 564640 495742
rect 564640 495662 564720 495742
rect 564720 495662 564748 495742
rect 564984 495662 565040 495742
rect 565040 495662 565120 495742
rect 565120 495662 565200 495742
rect 565200 495662 565220 495742
rect 565456 495662 565520 495742
rect 565520 495662 565600 495742
rect 565600 495662 565680 495742
rect 565680 495662 565692 495742
rect 565928 495662 566000 495742
rect 566000 495662 566080 495742
rect 566080 495662 566160 495742
rect 566160 495662 566164 495742
rect 566400 495662 566480 495742
rect 566480 495662 566560 495742
rect 566560 495662 566636 495742
rect 566872 495662 566880 495742
rect 566880 495662 566960 495742
rect 566960 495662 567040 495742
rect 567040 495662 567108 495742
rect 562624 495582 562860 495662
rect 563096 495582 563332 495662
rect 563568 495582 563804 495662
rect 564040 495582 564276 495662
rect 564512 495582 564748 495662
rect 564984 495582 565220 495662
rect 565456 495582 565692 495662
rect 565928 495582 566164 495662
rect 566400 495582 566636 495662
rect 566872 495582 567108 495662
rect 562624 495546 562640 495582
rect 562640 495546 562720 495582
rect 562720 495546 562800 495582
rect 562800 495546 562860 495582
rect 563096 495546 563120 495582
rect 563120 495546 563200 495582
rect 563200 495546 563280 495582
rect 563280 495546 563332 495582
rect 563568 495546 563600 495582
rect 563600 495546 563680 495582
rect 563680 495546 563760 495582
rect 563760 495546 563804 495582
rect 564040 495546 564080 495582
rect 564080 495546 564160 495582
rect 564160 495546 564240 495582
rect 564240 495546 564276 495582
rect 564512 495546 564560 495582
rect 564560 495546 564640 495582
rect 564640 495546 564720 495582
rect 564720 495546 564748 495582
rect 564984 495546 565040 495582
rect 565040 495546 565120 495582
rect 565120 495546 565200 495582
rect 565200 495546 565220 495582
rect 565456 495546 565520 495582
rect 565520 495546 565600 495582
rect 565600 495546 565680 495582
rect 565680 495546 565692 495582
rect 565928 495546 566000 495582
rect 566000 495546 566080 495582
rect 566080 495546 566160 495582
rect 566160 495546 566164 495582
rect 566400 495546 566480 495582
rect 566480 495546 566560 495582
rect 566560 495546 566636 495582
rect 566872 495546 566880 495582
rect 566880 495546 566960 495582
rect 566960 495546 567040 495582
rect 567040 495546 567108 495582
rect 572784 495742 573020 495782
rect 573256 495742 573492 495782
rect 573728 495742 573964 495782
rect 574200 495742 574436 495782
rect 574672 495742 574908 495782
rect 575144 495742 575380 495782
rect 575616 495742 575852 495782
rect 576088 495742 576324 495782
rect 576560 495742 576796 495782
rect 577032 495742 577268 495782
rect 572784 495662 572800 495742
rect 572800 495662 572880 495742
rect 572880 495662 572960 495742
rect 572960 495662 573020 495742
rect 573256 495662 573280 495742
rect 573280 495662 573360 495742
rect 573360 495662 573440 495742
rect 573440 495662 573492 495742
rect 573728 495662 573760 495742
rect 573760 495662 573840 495742
rect 573840 495662 573920 495742
rect 573920 495662 573964 495742
rect 574200 495662 574240 495742
rect 574240 495662 574320 495742
rect 574320 495662 574400 495742
rect 574400 495662 574436 495742
rect 574672 495662 574720 495742
rect 574720 495662 574800 495742
rect 574800 495662 574880 495742
rect 574880 495662 574908 495742
rect 575144 495662 575200 495742
rect 575200 495662 575280 495742
rect 575280 495662 575360 495742
rect 575360 495662 575380 495742
rect 575616 495662 575680 495742
rect 575680 495662 575760 495742
rect 575760 495662 575840 495742
rect 575840 495662 575852 495742
rect 576088 495662 576160 495742
rect 576160 495662 576240 495742
rect 576240 495662 576320 495742
rect 576320 495662 576324 495742
rect 576560 495662 576640 495742
rect 576640 495662 576720 495742
rect 576720 495662 576796 495742
rect 577032 495662 577040 495742
rect 577040 495662 577120 495742
rect 577120 495662 577200 495742
rect 577200 495662 577268 495742
rect 572784 495582 573020 495662
rect 573256 495582 573492 495662
rect 573728 495582 573964 495662
rect 574200 495582 574436 495662
rect 574672 495582 574908 495662
rect 575144 495582 575380 495662
rect 575616 495582 575852 495662
rect 576088 495582 576324 495662
rect 576560 495582 576796 495662
rect 577032 495582 577268 495662
rect 572784 495546 572800 495582
rect 572800 495546 572880 495582
rect 572880 495546 572960 495582
rect 572960 495546 573020 495582
rect 573256 495546 573280 495582
rect 573280 495546 573360 495582
rect 573360 495546 573440 495582
rect 573440 495546 573492 495582
rect 573728 495546 573760 495582
rect 573760 495546 573840 495582
rect 573840 495546 573920 495582
rect 573920 495546 573964 495582
rect 574200 495546 574240 495582
rect 574240 495546 574320 495582
rect 574320 495546 574400 495582
rect 574400 495546 574436 495582
rect 574672 495546 574720 495582
rect 574720 495546 574800 495582
rect 574800 495546 574880 495582
rect 574880 495546 574908 495582
rect 575144 495546 575200 495582
rect 575200 495546 575280 495582
rect 575280 495546 575360 495582
rect 575360 495546 575380 495582
rect 575616 495546 575680 495582
rect 575680 495546 575760 495582
rect 575760 495546 575840 495582
rect 575840 495546 575852 495582
rect 576088 495546 576160 495582
rect 576160 495546 576240 495582
rect 576240 495546 576320 495582
rect 576320 495546 576324 495582
rect 576560 495546 576640 495582
rect 576640 495546 576720 495582
rect 576720 495546 576796 495582
rect 577032 495546 577040 495582
rect 577040 495546 577120 495582
rect 577120 495546 577200 495582
rect 577200 495546 577268 495582
rect 572772 483800 573008 484036
rect 572772 483328 573008 483564
rect 572772 482856 573008 483092
rect 572772 482384 573008 482620
rect 572772 481912 573008 482148
rect 572772 481440 573008 481676
rect 572772 480968 573008 481204
rect 572772 480496 573008 480732
rect 572772 480024 573008 480260
rect 572772 479552 573008 479788
rect 572772 479080 573008 479316
rect 572772 478608 573008 478844
rect 572772 478136 573008 478372
rect 572772 477664 573008 477900
rect 573244 483800 573480 484036
rect 573244 483328 573480 483564
rect 573244 482856 573480 483092
rect 573244 482384 573480 482620
rect 573244 481912 573480 482148
rect 573244 481440 573480 481676
rect 573244 480968 573480 481204
rect 573244 480496 573480 480732
rect 573244 480024 573480 480260
rect 573244 479552 573480 479788
rect 573244 479080 573480 479316
rect 573244 478608 573480 478844
rect 573244 478136 573480 478372
rect 573244 477664 573480 477900
rect 573716 483800 573952 484036
rect 573716 483328 573952 483564
rect 573716 482856 573952 483092
rect 573716 482384 573952 482620
rect 573716 481912 573952 482148
rect 573716 481440 573952 481676
rect 573716 480968 573952 481204
rect 573716 480496 573952 480732
rect 573716 480024 573952 480260
rect 573716 479552 573952 479788
rect 573716 479080 573952 479316
rect 573716 478608 573952 478844
rect 573716 478136 573952 478372
rect 573716 477664 573952 477900
rect 574188 483800 574424 484036
rect 574188 483328 574424 483564
rect 574188 482856 574424 483092
rect 574188 482384 574424 482620
rect 574188 481912 574424 482148
rect 574188 481440 574424 481676
rect 574188 480968 574424 481204
rect 574188 480496 574424 480732
rect 574188 480024 574424 480260
rect 574188 479552 574424 479788
rect 574188 479080 574424 479316
rect 574188 478608 574424 478844
rect 574188 478136 574424 478372
rect 574188 477664 574424 477900
rect 574660 483800 574896 484036
rect 574660 483328 574896 483564
rect 574660 482856 574896 483092
rect 574660 482384 574896 482620
rect 574660 481912 574896 482148
rect 574660 481440 574896 481676
rect 574660 480968 574896 481204
rect 574660 480496 574896 480732
rect 574660 480024 574896 480260
rect 574660 479552 574896 479788
rect 574660 479080 574896 479316
rect 574660 478608 574896 478844
rect 574660 478136 574896 478372
rect 574660 477664 574896 477900
rect 575132 483800 575368 484036
rect 575132 483328 575368 483564
rect 575132 482856 575368 483092
rect 575132 482384 575368 482620
rect 575132 481912 575368 482148
rect 575132 481440 575368 481676
rect 575132 480968 575368 481204
rect 575132 480496 575368 480732
rect 575132 480024 575368 480260
rect 575132 479552 575368 479788
rect 575132 479080 575368 479316
rect 575132 478608 575368 478844
rect 575132 478136 575368 478372
rect 575132 477664 575368 477900
rect 575604 483800 575840 484036
rect 575604 483328 575840 483564
rect 575604 482856 575840 483092
rect 575604 482384 575840 482620
rect 575604 481912 575840 482148
rect 575604 481440 575840 481676
rect 575604 480968 575840 481204
rect 575604 480496 575840 480732
rect 575604 480024 575840 480260
rect 575604 479552 575840 479788
rect 575604 479080 575840 479316
rect 575604 478608 575840 478844
rect 575604 478136 575840 478372
rect 575604 477664 575840 477900
rect 576076 483800 576312 484036
rect 576076 483328 576312 483564
rect 576076 482856 576312 483092
rect 576076 482384 576312 482620
rect 576076 481912 576312 482148
rect 576076 481440 576312 481676
rect 576076 480968 576312 481204
rect 576076 480496 576312 480732
rect 576076 480024 576312 480260
rect 576076 479552 576312 479788
rect 576076 479080 576312 479316
rect 576076 478608 576312 478844
rect 576076 478136 576312 478372
rect 576076 477664 576312 477900
rect 576548 483800 576784 484036
rect 576548 483328 576784 483564
rect 576548 482856 576784 483092
rect 576548 482384 576784 482620
rect 576548 481912 576784 482148
rect 576548 481440 576784 481676
rect 576548 480968 576784 481204
rect 576548 480496 576784 480732
rect 576548 480024 576784 480260
rect 576548 479552 576784 479788
rect 576548 479080 576784 479316
rect 576548 478608 576784 478844
rect 576548 478136 576784 478372
rect 576548 477664 576784 477900
rect 577020 483800 577256 484036
rect 577020 483328 577256 483564
rect 577020 482856 577256 483092
rect 577020 482384 577256 482620
rect 577020 481912 577256 482148
rect 577020 481440 577256 481676
rect 577020 480968 577256 481204
rect 577020 480496 577256 480732
rect 577020 480024 577256 480260
rect 577020 479552 577256 479788
rect 577020 479080 577256 479316
rect 577020 478608 577256 478844
rect 577020 478136 577256 478372
rect 577020 477664 577256 477900
rect 512234 439888 513206 460198
rect 562624 455440 562860 455480
rect 563096 455440 563332 455480
rect 563568 455440 563804 455480
rect 564040 455440 564276 455480
rect 564512 455440 564748 455480
rect 564984 455440 565220 455480
rect 565456 455440 565692 455480
rect 565928 455440 566164 455480
rect 566400 455440 566636 455480
rect 566872 455440 567108 455480
rect 562624 455360 562640 455440
rect 562640 455360 562720 455440
rect 562720 455360 562800 455440
rect 562800 455360 562860 455440
rect 563096 455360 563120 455440
rect 563120 455360 563200 455440
rect 563200 455360 563280 455440
rect 563280 455360 563332 455440
rect 563568 455360 563600 455440
rect 563600 455360 563680 455440
rect 563680 455360 563760 455440
rect 563760 455360 563804 455440
rect 564040 455360 564080 455440
rect 564080 455360 564160 455440
rect 564160 455360 564240 455440
rect 564240 455360 564276 455440
rect 564512 455360 564560 455440
rect 564560 455360 564640 455440
rect 564640 455360 564720 455440
rect 564720 455360 564748 455440
rect 564984 455360 565040 455440
rect 565040 455360 565120 455440
rect 565120 455360 565200 455440
rect 565200 455360 565220 455440
rect 565456 455360 565520 455440
rect 565520 455360 565600 455440
rect 565600 455360 565680 455440
rect 565680 455360 565692 455440
rect 565928 455360 566000 455440
rect 566000 455360 566080 455440
rect 566080 455360 566160 455440
rect 566160 455360 566164 455440
rect 566400 455360 566480 455440
rect 566480 455360 566560 455440
rect 566560 455360 566636 455440
rect 566872 455360 566880 455440
rect 566880 455360 566960 455440
rect 566960 455360 567040 455440
rect 567040 455360 567108 455440
rect 562624 455280 562860 455360
rect 563096 455280 563332 455360
rect 563568 455280 563804 455360
rect 564040 455280 564276 455360
rect 564512 455280 564748 455360
rect 564984 455280 565220 455360
rect 565456 455280 565692 455360
rect 565928 455280 566164 455360
rect 566400 455280 566636 455360
rect 566872 455280 567108 455360
rect 562624 455244 562640 455280
rect 562640 455244 562720 455280
rect 562720 455244 562800 455280
rect 562800 455244 562860 455280
rect 563096 455244 563120 455280
rect 563120 455244 563200 455280
rect 563200 455244 563280 455280
rect 563280 455244 563332 455280
rect 563568 455244 563600 455280
rect 563600 455244 563680 455280
rect 563680 455244 563760 455280
rect 563760 455244 563804 455280
rect 564040 455244 564080 455280
rect 564080 455244 564160 455280
rect 564160 455244 564240 455280
rect 564240 455244 564276 455280
rect 564512 455244 564560 455280
rect 564560 455244 564640 455280
rect 564640 455244 564720 455280
rect 564720 455244 564748 455280
rect 564984 455244 565040 455280
rect 565040 455244 565120 455280
rect 565120 455244 565200 455280
rect 565200 455244 565220 455280
rect 565456 455244 565520 455280
rect 565520 455244 565600 455280
rect 565600 455244 565680 455280
rect 565680 455244 565692 455280
rect 565928 455244 566000 455280
rect 566000 455244 566080 455280
rect 566080 455244 566160 455280
rect 566160 455244 566164 455280
rect 566400 455244 566480 455280
rect 566480 455244 566560 455280
rect 566560 455244 566636 455280
rect 566872 455244 566880 455280
rect 566880 455244 566960 455280
rect 566960 455244 567040 455280
rect 567040 455244 567108 455280
rect 572784 455440 573020 455480
rect 573256 455440 573492 455480
rect 573728 455440 573964 455480
rect 574200 455440 574436 455480
rect 574672 455440 574908 455480
rect 575144 455440 575380 455480
rect 575616 455440 575852 455480
rect 576088 455440 576324 455480
rect 576560 455440 576796 455480
rect 577032 455440 577268 455480
rect 572784 455360 572800 455440
rect 572800 455360 572880 455440
rect 572880 455360 572960 455440
rect 572960 455360 573020 455440
rect 573256 455360 573280 455440
rect 573280 455360 573360 455440
rect 573360 455360 573440 455440
rect 573440 455360 573492 455440
rect 573728 455360 573760 455440
rect 573760 455360 573840 455440
rect 573840 455360 573920 455440
rect 573920 455360 573964 455440
rect 574200 455360 574240 455440
rect 574240 455360 574320 455440
rect 574320 455360 574400 455440
rect 574400 455360 574436 455440
rect 574672 455360 574720 455440
rect 574720 455360 574800 455440
rect 574800 455360 574880 455440
rect 574880 455360 574908 455440
rect 575144 455360 575200 455440
rect 575200 455360 575280 455440
rect 575280 455360 575360 455440
rect 575360 455360 575380 455440
rect 575616 455360 575680 455440
rect 575680 455360 575760 455440
rect 575760 455360 575840 455440
rect 575840 455360 575852 455440
rect 576088 455360 576160 455440
rect 576160 455360 576240 455440
rect 576240 455360 576320 455440
rect 576320 455360 576324 455440
rect 576560 455360 576640 455440
rect 576640 455360 576720 455440
rect 576720 455360 576796 455440
rect 577032 455360 577040 455440
rect 577040 455360 577120 455440
rect 577120 455360 577200 455440
rect 577200 455360 577268 455440
rect 572784 455280 573020 455360
rect 573256 455280 573492 455360
rect 573728 455280 573964 455360
rect 574200 455280 574436 455360
rect 574672 455280 574908 455360
rect 575144 455280 575380 455360
rect 575616 455280 575852 455360
rect 576088 455280 576324 455360
rect 576560 455280 576796 455360
rect 577032 455280 577268 455360
rect 572784 455244 572800 455280
rect 572800 455244 572880 455280
rect 572880 455244 572960 455280
rect 572960 455244 573020 455280
rect 573256 455244 573280 455280
rect 573280 455244 573360 455280
rect 573360 455244 573440 455280
rect 573440 455244 573492 455280
rect 573728 455244 573760 455280
rect 573760 455244 573840 455280
rect 573840 455244 573920 455280
rect 573920 455244 573964 455280
rect 574200 455244 574240 455280
rect 574240 455244 574320 455280
rect 574320 455244 574400 455280
rect 574400 455244 574436 455280
rect 574672 455244 574720 455280
rect 574720 455244 574800 455280
rect 574800 455244 574880 455280
rect 574880 455244 574908 455280
rect 575144 455244 575200 455280
rect 575200 455244 575280 455280
rect 575280 455244 575360 455280
rect 575360 455244 575380 455280
rect 575616 455244 575680 455280
rect 575680 455244 575760 455280
rect 575760 455244 575840 455280
rect 575840 455244 575852 455280
rect 576088 455244 576160 455280
rect 576160 455244 576240 455280
rect 576240 455244 576320 455280
rect 576320 455244 576324 455280
rect 576560 455244 576640 455280
rect 576640 455244 576720 455280
rect 576720 455244 576796 455280
rect 577032 455244 577040 455280
rect 577040 455244 577120 455280
rect 577120 455244 577200 455280
rect 577200 455244 577268 455280
rect 572772 426452 573008 426688
rect 572772 425980 573008 426216
rect 572772 425508 573008 425744
rect 572772 425036 573008 425272
rect 572772 424564 573008 424800
rect 572772 424092 573008 424328
rect 572772 423620 573008 423856
rect 572772 423148 573008 423384
rect 572772 422676 573008 422912
rect 572772 422204 573008 422440
rect 572772 421732 573008 421968
rect 572772 421260 573008 421496
rect 572772 420788 573008 421024
rect 572772 420316 573008 420552
rect 573244 426452 573480 426688
rect 573244 425980 573480 426216
rect 573244 425508 573480 425744
rect 573244 425036 573480 425272
rect 573244 424564 573480 424800
rect 573244 424092 573480 424328
rect 573244 423620 573480 423856
rect 573244 423148 573480 423384
rect 573244 422676 573480 422912
rect 573244 422204 573480 422440
rect 573244 421732 573480 421968
rect 573244 421260 573480 421496
rect 573244 420788 573480 421024
rect 573244 420316 573480 420552
rect 573716 426452 573952 426688
rect 573716 425980 573952 426216
rect 573716 425508 573952 425744
rect 573716 425036 573952 425272
rect 573716 424564 573952 424800
rect 573716 424092 573952 424328
rect 573716 423620 573952 423856
rect 573716 423148 573952 423384
rect 573716 422676 573952 422912
rect 573716 422204 573952 422440
rect 573716 421732 573952 421968
rect 573716 421260 573952 421496
rect 573716 420788 573952 421024
rect 573716 420316 573952 420552
rect 574188 426452 574424 426688
rect 574188 425980 574424 426216
rect 574188 425508 574424 425744
rect 574188 425036 574424 425272
rect 574188 424564 574424 424800
rect 574188 424092 574424 424328
rect 574188 423620 574424 423856
rect 574188 423148 574424 423384
rect 574188 422676 574424 422912
rect 574188 422204 574424 422440
rect 574188 421732 574424 421968
rect 574188 421260 574424 421496
rect 574188 420788 574424 421024
rect 574188 420316 574424 420552
rect 574660 426452 574896 426688
rect 574660 425980 574896 426216
rect 574660 425508 574896 425744
rect 574660 425036 574896 425272
rect 574660 424564 574896 424800
rect 574660 424092 574896 424328
rect 574660 423620 574896 423856
rect 574660 423148 574896 423384
rect 574660 422676 574896 422912
rect 574660 422204 574896 422440
rect 574660 421732 574896 421968
rect 574660 421260 574896 421496
rect 574660 420788 574896 421024
rect 574660 420316 574896 420552
rect 575132 426452 575368 426688
rect 575132 425980 575368 426216
rect 575132 425508 575368 425744
rect 575132 425036 575368 425272
rect 575132 424564 575368 424800
rect 575132 424092 575368 424328
rect 575132 423620 575368 423856
rect 575132 423148 575368 423384
rect 575132 422676 575368 422912
rect 575132 422204 575368 422440
rect 575132 421732 575368 421968
rect 575132 421260 575368 421496
rect 575132 420788 575368 421024
rect 575132 420316 575368 420552
rect 575604 426452 575840 426688
rect 575604 425980 575840 426216
rect 575604 425508 575840 425744
rect 575604 425036 575840 425272
rect 575604 424564 575840 424800
rect 575604 424092 575840 424328
rect 575604 423620 575840 423856
rect 575604 423148 575840 423384
rect 575604 422676 575840 422912
rect 575604 422204 575840 422440
rect 575604 421732 575840 421968
rect 575604 421260 575840 421496
rect 575604 420788 575840 421024
rect 575604 420316 575840 420552
rect 576076 426452 576312 426688
rect 576076 425980 576312 426216
rect 576076 425508 576312 425744
rect 576076 425036 576312 425272
rect 576076 424564 576312 424800
rect 576076 424092 576312 424328
rect 576076 423620 576312 423856
rect 576076 423148 576312 423384
rect 576076 422676 576312 422912
rect 576076 422204 576312 422440
rect 576076 421732 576312 421968
rect 576076 421260 576312 421496
rect 576076 420788 576312 421024
rect 576076 420316 576312 420552
rect 576548 426452 576784 426688
rect 576548 425980 576784 426216
rect 576548 425508 576784 425744
rect 576548 425036 576784 425272
rect 576548 424564 576784 424800
rect 576548 424092 576784 424328
rect 576548 423620 576784 423856
rect 576548 423148 576784 423384
rect 576548 422676 576784 422912
rect 576548 422204 576784 422440
rect 576548 421732 576784 421968
rect 576548 421260 576784 421496
rect 576548 420788 576784 421024
rect 576548 420316 576784 420552
rect 577020 426452 577256 426688
rect 577020 425980 577256 426216
rect 577020 425508 577256 425744
rect 577020 425036 577256 425272
rect 577020 424564 577256 424800
rect 577020 424092 577256 424328
rect 577020 423620 577256 423856
rect 577020 423148 577256 423384
rect 577020 422676 577256 422912
rect 577020 422204 577256 422440
rect 577020 421732 577256 421968
rect 577020 421260 577256 421496
rect 577020 420788 577256 421024
rect 577020 420316 577256 420552
rect 562624 377128 562860 377364
rect 562624 376656 562860 376892
rect 562624 376184 562860 376420
rect 562624 375712 562860 375948
rect 562624 375240 562860 375476
rect 562624 374768 562860 375004
rect 562624 374296 562860 374532
rect 562624 373824 562860 374060
rect 562624 373352 562860 373588
rect 562624 372880 562860 373116
rect 562624 372408 562860 372644
rect 562624 371936 562860 372172
rect 562624 371464 562860 371700
rect 563096 377128 563332 377364
rect 563096 376656 563332 376892
rect 563096 376184 563332 376420
rect 563096 375712 563332 375948
rect 563096 375240 563332 375476
rect 563096 374768 563332 375004
rect 563096 374296 563332 374532
rect 563096 373824 563332 374060
rect 563096 373352 563332 373588
rect 563096 372880 563332 373116
rect 563096 372408 563332 372644
rect 563096 371936 563332 372172
rect 563096 371464 563332 371700
rect 563568 377128 563804 377364
rect 563568 376656 563804 376892
rect 563568 376184 563804 376420
rect 563568 375712 563804 375948
rect 563568 375240 563804 375476
rect 563568 374768 563804 375004
rect 563568 374296 563804 374532
rect 563568 373824 563804 374060
rect 563568 373352 563804 373588
rect 563568 372880 563804 373116
rect 563568 372408 563804 372644
rect 563568 371936 563804 372172
rect 563568 371464 563804 371700
rect 564040 377128 564276 377364
rect 564040 376656 564276 376892
rect 564040 376184 564276 376420
rect 564040 375712 564276 375948
rect 564040 375240 564276 375476
rect 564040 374768 564276 375004
rect 564040 374296 564276 374532
rect 564040 373824 564276 374060
rect 564040 373352 564276 373588
rect 564040 372880 564276 373116
rect 564040 372408 564276 372644
rect 564040 371936 564276 372172
rect 564040 371464 564276 371700
rect 564512 377128 564748 377364
rect 564512 376656 564748 376892
rect 564512 376184 564748 376420
rect 564512 375712 564748 375948
rect 564512 375240 564748 375476
rect 564512 374768 564748 375004
rect 564512 374296 564748 374532
rect 564512 373824 564748 374060
rect 564512 373352 564748 373588
rect 564512 372880 564748 373116
rect 564512 372408 564748 372644
rect 564512 371936 564748 372172
rect 564512 371464 564748 371700
rect 564984 377128 565220 377364
rect 564984 376656 565220 376892
rect 564984 376184 565220 376420
rect 564984 375712 565220 375948
rect 564984 375240 565220 375476
rect 564984 374768 565220 375004
rect 564984 374296 565220 374532
rect 564984 373824 565220 374060
rect 564984 373352 565220 373588
rect 564984 372880 565220 373116
rect 564984 372408 565220 372644
rect 564984 371936 565220 372172
rect 564984 371464 565220 371700
rect 565456 377128 565692 377364
rect 565456 376656 565692 376892
rect 565456 376184 565692 376420
rect 565456 375712 565692 375948
rect 565456 375240 565692 375476
rect 565456 374768 565692 375004
rect 565456 374296 565692 374532
rect 565456 373824 565692 374060
rect 565456 373352 565692 373588
rect 565456 372880 565692 373116
rect 565456 372408 565692 372644
rect 565456 371936 565692 372172
rect 565456 371464 565692 371700
rect 565928 377128 566164 377364
rect 565928 376656 566164 376892
rect 565928 376184 566164 376420
rect 565928 375712 566164 375948
rect 565928 375240 566164 375476
rect 565928 374768 566164 375004
rect 565928 374296 566164 374532
rect 565928 373824 566164 374060
rect 565928 373352 566164 373588
rect 565928 372880 566164 373116
rect 565928 372408 566164 372644
rect 565928 371936 566164 372172
rect 565928 371464 566164 371700
rect 566400 377128 566636 377364
rect 566400 376656 566636 376892
rect 566400 376184 566636 376420
rect 566400 375712 566636 375948
rect 566400 375240 566636 375476
rect 566400 374768 566636 375004
rect 566400 374296 566636 374532
rect 566400 373824 566636 374060
rect 566400 373352 566636 373588
rect 566400 372880 566636 373116
rect 566400 372408 566636 372644
rect 566400 371936 566636 372172
rect 566400 371464 566636 371700
rect 566872 377128 567108 377364
rect 566872 376656 567108 376892
rect 566872 376184 567108 376420
rect 566872 375712 567108 375948
rect 566872 375240 567108 375476
rect 566872 374768 567108 375004
rect 566872 374296 567108 374532
rect 566872 373824 567108 374060
rect 566872 373352 567108 373588
rect 566872 372880 567108 373116
rect 566872 372408 567108 372644
rect 566872 371936 567108 372172
rect 566872 371464 567108 371700
<< mimcap2 >>
rect 518532 472390 518932 472430
rect 518532 472070 518572 472390
rect 518892 472070 518932 472390
rect 518532 472030 518932 472070
rect 519232 472390 519632 472430
rect 519232 472070 519272 472390
rect 519592 472070 519632 472390
rect 519232 472030 519632 472070
rect 519932 472390 520332 472430
rect 519932 472070 519972 472390
rect 520292 472070 520332 472390
rect 519932 472030 520332 472070
rect 520632 472390 521032 472430
rect 520632 472070 520672 472390
rect 520992 472070 521032 472390
rect 520632 472030 521032 472070
rect 521332 472390 521732 472430
rect 521332 472070 521372 472390
rect 521692 472070 521732 472390
rect 521332 472030 521732 472070
rect 522032 472390 522432 472430
rect 522032 472070 522072 472390
rect 522392 472070 522432 472390
rect 522032 472030 522432 472070
rect 522732 472390 523132 472430
rect 522732 472070 522772 472390
rect 523092 472070 523132 472390
rect 522732 472030 523132 472070
rect 523432 472390 523832 472430
rect 523432 472070 523472 472390
rect 523792 472070 523832 472390
rect 523432 472030 523832 472070
rect 524132 472390 524532 472430
rect 524132 472070 524172 472390
rect 524492 472070 524532 472390
rect 524132 472030 524532 472070
rect 524832 472390 525232 472430
rect 524832 472070 524872 472390
rect 525192 472070 525232 472390
rect 524832 472030 525232 472070
rect 518532 471268 518932 471308
rect 518532 470948 518572 471268
rect 518892 470948 518932 471268
rect 518532 470908 518932 470948
rect 519232 471268 519632 471308
rect 519232 470948 519272 471268
rect 519592 470948 519632 471268
rect 519232 470908 519632 470948
rect 519932 471268 520332 471308
rect 519932 470948 519972 471268
rect 520292 470948 520332 471268
rect 519932 470908 520332 470948
rect 520632 471268 521032 471308
rect 520632 470948 520672 471268
rect 520992 470948 521032 471268
rect 520632 470908 521032 470948
rect 521332 471268 521732 471308
rect 521332 470948 521372 471268
rect 521692 470948 521732 471268
rect 521332 470908 521732 470948
rect 522032 471268 522432 471308
rect 522032 470948 522072 471268
rect 522392 470948 522432 471268
rect 522032 470908 522432 470948
rect 522732 471268 523132 471308
rect 522732 470948 522772 471268
rect 523092 470948 523132 471268
rect 522732 470908 523132 470948
rect 523432 471268 523832 471308
rect 523432 470948 523472 471268
rect 523792 470948 523832 471268
rect 523432 470908 523832 470948
rect 524132 471268 524532 471308
rect 524132 470948 524172 471268
rect 524492 470948 524532 471268
rect 524132 470908 524532 470948
rect 524832 471268 525232 471308
rect 524832 470948 524872 471268
rect 525192 470948 525232 471268
rect 524832 470908 525232 470948
rect 518532 470146 518932 470186
rect 518532 469826 518572 470146
rect 518892 469826 518932 470146
rect 518532 469786 518932 469826
rect 519232 470146 519632 470186
rect 519232 469826 519272 470146
rect 519592 469826 519632 470146
rect 519232 469786 519632 469826
rect 519932 470146 520332 470186
rect 519932 469826 519972 470146
rect 520292 469826 520332 470146
rect 519932 469786 520332 469826
rect 520632 470146 521032 470186
rect 520632 469826 520672 470146
rect 520992 469826 521032 470146
rect 520632 469786 521032 469826
rect 521332 470146 521732 470186
rect 521332 469826 521372 470146
rect 521692 469826 521732 470146
rect 521332 469786 521732 469826
rect 522032 470146 522432 470186
rect 522032 469826 522072 470146
rect 522392 469826 522432 470146
rect 522032 469786 522432 469826
rect 522732 470146 523132 470186
rect 522732 469826 522772 470146
rect 523092 469826 523132 470146
rect 522732 469786 523132 469826
rect 523432 470146 523832 470186
rect 523432 469826 523472 470146
rect 523792 469826 523832 470146
rect 523432 469786 523832 469826
rect 524132 470146 524532 470186
rect 524132 469826 524172 470146
rect 524492 469826 524532 470146
rect 524132 469786 524532 469826
rect 524832 470146 525232 470186
rect 524832 469826 524872 470146
rect 525192 469826 525232 470146
rect 524832 469786 525232 469826
rect 518532 469024 518932 469064
rect 518532 468704 518572 469024
rect 518892 468704 518932 469024
rect 518532 468664 518932 468704
rect 519232 469024 519632 469064
rect 519232 468704 519272 469024
rect 519592 468704 519632 469024
rect 519232 468664 519632 468704
rect 519932 469024 520332 469064
rect 519932 468704 519972 469024
rect 520292 468704 520332 469024
rect 519932 468664 520332 468704
rect 520632 469024 521032 469064
rect 520632 468704 520672 469024
rect 520992 468704 521032 469024
rect 520632 468664 521032 468704
rect 521332 469024 521732 469064
rect 521332 468704 521372 469024
rect 521692 468704 521732 469024
rect 521332 468664 521732 468704
rect 522032 469024 522432 469064
rect 522032 468704 522072 469024
rect 522392 468704 522432 469024
rect 522032 468664 522432 468704
rect 522732 469024 523132 469064
rect 522732 468704 522772 469024
rect 523092 468704 523132 469024
rect 522732 468664 523132 468704
rect 523432 469024 523832 469064
rect 523432 468704 523472 469024
rect 523792 468704 523832 469024
rect 523432 468664 523832 468704
rect 524132 469024 524532 469064
rect 524132 468704 524172 469024
rect 524492 468704 524532 469024
rect 524132 468664 524532 468704
rect 524832 469024 525232 469064
rect 524832 468704 524872 469024
rect 525192 468704 525232 469024
rect 524832 468664 525232 468704
rect 518532 467902 518932 467942
rect 518532 467582 518572 467902
rect 518892 467582 518932 467902
rect 518532 467542 518932 467582
rect 519232 467902 519632 467942
rect 519232 467582 519272 467902
rect 519592 467582 519632 467902
rect 519232 467542 519632 467582
rect 519932 467902 520332 467942
rect 519932 467582 519972 467902
rect 520292 467582 520332 467902
rect 519932 467542 520332 467582
rect 520632 467902 521032 467942
rect 520632 467582 520672 467902
rect 520992 467582 521032 467902
rect 520632 467542 521032 467582
rect 521332 467902 521732 467942
rect 521332 467582 521372 467902
rect 521692 467582 521732 467902
rect 521332 467542 521732 467582
rect 522032 467902 522432 467942
rect 522032 467582 522072 467902
rect 522392 467582 522432 467902
rect 522032 467542 522432 467582
rect 522732 467902 523132 467942
rect 522732 467582 522772 467902
rect 523092 467582 523132 467902
rect 522732 467542 523132 467582
rect 523432 467902 523832 467942
rect 523432 467582 523472 467902
rect 523792 467582 523832 467902
rect 523432 467542 523832 467582
rect 524132 467902 524532 467942
rect 524132 467582 524172 467902
rect 524492 467582 524532 467902
rect 524132 467542 524532 467582
rect 524832 467902 525232 467942
rect 524832 467582 524872 467902
rect 525192 467582 525232 467902
rect 524832 467542 525232 467582
rect 518532 466780 518932 466820
rect 518532 466460 518572 466780
rect 518892 466460 518932 466780
rect 518532 466420 518932 466460
rect 519232 466780 519632 466820
rect 519232 466460 519272 466780
rect 519592 466460 519632 466780
rect 519232 466420 519632 466460
rect 519932 466780 520332 466820
rect 519932 466460 519972 466780
rect 520292 466460 520332 466780
rect 519932 466420 520332 466460
rect 520632 466780 521032 466820
rect 520632 466460 520672 466780
rect 520992 466460 521032 466780
rect 520632 466420 521032 466460
rect 521332 466780 521732 466820
rect 521332 466460 521372 466780
rect 521692 466460 521732 466780
rect 521332 466420 521732 466460
rect 522032 466780 522432 466820
rect 522032 466460 522072 466780
rect 522392 466460 522432 466780
rect 522032 466420 522432 466460
rect 522732 466780 523132 466820
rect 522732 466460 522772 466780
rect 523092 466460 523132 466780
rect 522732 466420 523132 466460
rect 523432 466780 523832 466820
rect 523432 466460 523472 466780
rect 523792 466460 523832 466780
rect 523432 466420 523832 466460
rect 524132 466780 524532 466820
rect 524132 466460 524172 466780
rect 524492 466460 524532 466780
rect 524132 466420 524532 466460
rect 524832 466780 525232 466820
rect 524832 466460 524872 466780
rect 525192 466460 525232 466780
rect 524832 466420 525232 466460
rect 518532 465658 518932 465698
rect 518532 465338 518572 465658
rect 518892 465338 518932 465658
rect 518532 465298 518932 465338
rect 519232 465658 519632 465698
rect 519232 465338 519272 465658
rect 519592 465338 519632 465658
rect 519232 465298 519632 465338
rect 519932 465658 520332 465698
rect 519932 465338 519972 465658
rect 520292 465338 520332 465658
rect 519932 465298 520332 465338
rect 520632 465658 521032 465698
rect 520632 465338 520672 465658
rect 520992 465338 521032 465658
rect 520632 465298 521032 465338
rect 521332 465658 521732 465698
rect 521332 465338 521372 465658
rect 521692 465338 521732 465658
rect 521332 465298 521732 465338
rect 522032 465658 522432 465698
rect 522032 465338 522072 465658
rect 522392 465338 522432 465658
rect 522032 465298 522432 465338
rect 522732 465658 523132 465698
rect 522732 465338 522772 465658
rect 523092 465338 523132 465658
rect 522732 465298 523132 465338
rect 523432 465658 523832 465698
rect 523432 465338 523472 465658
rect 523792 465338 523832 465658
rect 523432 465298 523832 465338
rect 524132 465658 524532 465698
rect 524132 465338 524172 465658
rect 524492 465338 524532 465658
rect 524132 465298 524532 465338
rect 524832 465658 525232 465698
rect 524832 465338 524872 465658
rect 525192 465338 525232 465658
rect 524832 465298 525232 465338
rect 518532 464536 518932 464576
rect 518532 464216 518572 464536
rect 518892 464216 518932 464536
rect 518532 464176 518932 464216
rect 519232 464536 519632 464576
rect 519232 464216 519272 464536
rect 519592 464216 519632 464536
rect 519232 464176 519632 464216
rect 519932 464536 520332 464576
rect 519932 464216 519972 464536
rect 520292 464216 520332 464536
rect 519932 464176 520332 464216
rect 520632 464536 521032 464576
rect 520632 464216 520672 464536
rect 520992 464216 521032 464536
rect 520632 464176 521032 464216
rect 521332 464536 521732 464576
rect 521332 464216 521372 464536
rect 521692 464216 521732 464536
rect 521332 464176 521732 464216
rect 522032 464536 522432 464576
rect 522032 464216 522072 464536
rect 522392 464216 522432 464536
rect 522032 464176 522432 464216
rect 522732 464536 523132 464576
rect 522732 464216 522772 464536
rect 523092 464216 523132 464536
rect 522732 464176 523132 464216
rect 523432 464536 523832 464576
rect 523432 464216 523472 464536
rect 523792 464216 523832 464536
rect 523432 464176 523832 464216
rect 524132 464536 524532 464576
rect 524132 464216 524172 464536
rect 524492 464216 524532 464536
rect 524132 464176 524532 464216
rect 524832 464536 525232 464576
rect 524832 464216 524872 464536
rect 525192 464216 525232 464536
rect 524832 464176 525232 464216
rect 518532 463414 518932 463454
rect 518532 463094 518572 463414
rect 518892 463094 518932 463414
rect 518532 463054 518932 463094
rect 519232 463414 519632 463454
rect 519232 463094 519272 463414
rect 519592 463094 519632 463414
rect 519232 463054 519632 463094
rect 519932 463414 520332 463454
rect 519932 463094 519972 463414
rect 520292 463094 520332 463414
rect 519932 463054 520332 463094
rect 520632 463414 521032 463454
rect 520632 463094 520672 463414
rect 520992 463094 521032 463414
rect 520632 463054 521032 463094
rect 521332 463414 521732 463454
rect 521332 463094 521372 463414
rect 521692 463094 521732 463414
rect 521332 463054 521732 463094
rect 522032 463414 522432 463454
rect 522032 463094 522072 463414
rect 522392 463094 522432 463414
rect 522032 463054 522432 463094
rect 522732 463414 523132 463454
rect 522732 463094 522772 463414
rect 523092 463094 523132 463414
rect 522732 463054 523132 463094
rect 523432 463414 523832 463454
rect 523432 463094 523472 463414
rect 523792 463094 523832 463414
rect 523432 463054 523832 463094
rect 524132 463414 524532 463454
rect 524132 463094 524172 463414
rect 524492 463094 524532 463414
rect 524132 463054 524532 463094
rect 524832 463414 525232 463454
rect 524832 463094 524872 463414
rect 525192 463094 525232 463414
rect 524832 463054 525232 463094
rect 518532 462292 518932 462332
rect 518532 461972 518572 462292
rect 518892 461972 518932 462292
rect 518532 461932 518932 461972
rect 519232 462292 519632 462332
rect 519232 461972 519272 462292
rect 519592 461972 519632 462292
rect 519232 461932 519632 461972
rect 519932 462292 520332 462332
rect 519932 461972 519972 462292
rect 520292 461972 520332 462292
rect 519932 461932 520332 461972
rect 520632 462292 521032 462332
rect 520632 461972 520672 462292
rect 520992 461972 521032 462292
rect 520632 461932 521032 461972
rect 521332 462292 521732 462332
rect 521332 461972 521372 462292
rect 521692 461972 521732 462292
rect 521332 461932 521732 461972
rect 522032 462292 522432 462332
rect 522032 461972 522072 462292
rect 522392 461972 522432 462292
rect 522032 461932 522432 461972
rect 522732 462292 523132 462332
rect 522732 461972 522772 462292
rect 523092 461972 523132 462292
rect 522732 461932 523132 461972
rect 523432 462292 523832 462332
rect 523432 461972 523472 462292
rect 523792 461972 523832 462292
rect 523432 461932 523832 461972
rect 524132 462292 524532 462332
rect 524132 461972 524172 462292
rect 524492 461972 524532 462292
rect 524132 461932 524532 461972
rect 524832 462292 525232 462332
rect 524832 461972 524872 462292
rect 525192 461972 525232 462292
rect 524832 461932 525232 461972
<< mimcap2contact >>
rect 518572 472070 518892 472390
rect 519272 472070 519592 472390
rect 519972 472070 520292 472390
rect 520672 472070 520992 472390
rect 521372 472070 521692 472390
rect 522072 472070 522392 472390
rect 522772 472070 523092 472390
rect 523472 472070 523792 472390
rect 524172 472070 524492 472390
rect 524872 472070 525192 472390
rect 518572 470948 518892 471268
rect 519272 470948 519592 471268
rect 519972 470948 520292 471268
rect 520672 470948 520992 471268
rect 521372 470948 521692 471268
rect 522072 470948 522392 471268
rect 522772 470948 523092 471268
rect 523472 470948 523792 471268
rect 524172 470948 524492 471268
rect 524872 470948 525192 471268
rect 518572 469826 518892 470146
rect 519272 469826 519592 470146
rect 519972 469826 520292 470146
rect 520672 469826 520992 470146
rect 521372 469826 521692 470146
rect 522072 469826 522392 470146
rect 522772 469826 523092 470146
rect 523472 469826 523792 470146
rect 524172 469826 524492 470146
rect 524872 469826 525192 470146
rect 518572 468704 518892 469024
rect 519272 468704 519592 469024
rect 519972 468704 520292 469024
rect 520672 468704 520992 469024
rect 521372 468704 521692 469024
rect 522072 468704 522392 469024
rect 522772 468704 523092 469024
rect 523472 468704 523792 469024
rect 524172 468704 524492 469024
rect 524872 468704 525192 469024
rect 518572 467582 518892 467902
rect 519272 467582 519592 467902
rect 519972 467582 520292 467902
rect 520672 467582 520992 467902
rect 521372 467582 521692 467902
rect 522072 467582 522392 467902
rect 522772 467582 523092 467902
rect 523472 467582 523792 467902
rect 524172 467582 524492 467902
rect 524872 467582 525192 467902
rect 518572 466460 518892 466780
rect 519272 466460 519592 466780
rect 519972 466460 520292 466780
rect 520672 466460 520992 466780
rect 521372 466460 521692 466780
rect 522072 466460 522392 466780
rect 522772 466460 523092 466780
rect 523472 466460 523792 466780
rect 524172 466460 524492 466780
rect 524872 466460 525192 466780
rect 518572 465338 518892 465658
rect 519272 465338 519592 465658
rect 519972 465338 520292 465658
rect 520672 465338 520992 465658
rect 521372 465338 521692 465658
rect 522072 465338 522392 465658
rect 522772 465338 523092 465658
rect 523472 465338 523792 465658
rect 524172 465338 524492 465658
rect 524872 465338 525192 465658
rect 518572 464216 518892 464536
rect 519272 464216 519592 464536
rect 519972 464216 520292 464536
rect 520672 464216 520992 464536
rect 521372 464216 521692 464536
rect 522072 464216 522392 464536
rect 522772 464216 523092 464536
rect 523472 464216 523792 464536
rect 524172 464216 524492 464536
rect 524872 464216 525192 464536
rect 518572 463094 518892 463414
rect 519272 463094 519592 463414
rect 519972 463094 520292 463414
rect 520672 463094 520992 463414
rect 521372 463094 521692 463414
rect 522072 463094 522392 463414
rect 522772 463094 523092 463414
rect 523472 463094 523792 463414
rect 524172 463094 524492 463414
rect 524872 463094 525192 463414
rect 518572 461972 518892 462292
rect 519272 461972 519592 462292
rect 519972 461972 520292 462292
rect 520672 461972 520992 462292
rect 521372 461972 521692 462292
rect 522072 461972 522392 462292
rect 522772 461972 523092 462292
rect 523472 461972 523792 462292
rect 524172 461972 524492 462292
rect 524872 461972 525192 462292
<< metal5 >>
rect 572560 697380 577480 697420
rect 572560 697144 577492 697380
rect 572560 696908 572772 697144
rect 573008 696908 573244 697144
rect 573480 696908 573716 697144
rect 573952 696908 574188 697144
rect 574424 696908 574660 697144
rect 574896 696908 575132 697144
rect 575368 696908 575604 697144
rect 575840 696908 576076 697144
rect 576312 696908 576548 697144
rect 576784 696908 577020 697144
rect 577256 696908 577492 697144
rect 572560 696672 577492 696908
rect 572560 696436 572772 696672
rect 573008 696436 573244 696672
rect 573480 696436 573716 696672
rect 573952 696436 574188 696672
rect 574424 696436 574660 696672
rect 574896 696436 575132 696672
rect 575368 696436 575604 696672
rect 575840 696436 576076 696672
rect 576312 696436 576548 696672
rect 576784 696436 577020 696672
rect 577256 696436 577492 696672
rect 572560 696200 577492 696436
rect 572560 695964 572772 696200
rect 573008 695964 573244 696200
rect 573480 695964 573716 696200
rect 573952 695964 574188 696200
rect 574424 695964 574660 696200
rect 574896 695964 575132 696200
rect 575368 695964 575604 696200
rect 575840 695964 576076 696200
rect 576312 695964 576548 696200
rect 576784 695964 577020 696200
rect 577256 695964 577492 696200
rect 572560 695728 577492 695964
rect 572560 695492 572772 695728
rect 573008 695492 573244 695728
rect 573480 695492 573716 695728
rect 573952 695492 574188 695728
rect 574424 695492 574660 695728
rect 574896 695492 575132 695728
rect 575368 695492 575604 695728
rect 575840 695492 576076 695728
rect 576312 695492 576548 695728
rect 576784 695492 577020 695728
rect 577256 695492 577492 695728
rect 572560 695256 577492 695492
rect 572560 695020 572772 695256
rect 573008 695020 573244 695256
rect 573480 695020 573716 695256
rect 573952 695020 574188 695256
rect 574424 695020 574660 695256
rect 574896 695020 575132 695256
rect 575368 695020 575604 695256
rect 575840 695020 576076 695256
rect 576312 695020 576548 695256
rect 576784 695020 577020 695256
rect 577256 695020 577492 695256
rect 572560 694784 577492 695020
rect 572560 694548 572772 694784
rect 573008 694548 573244 694784
rect 573480 694548 573716 694784
rect 573952 694548 574188 694784
rect 574424 694548 574660 694784
rect 574896 694548 575132 694784
rect 575368 694548 575604 694784
rect 575840 694548 576076 694784
rect 576312 694548 576548 694784
rect 576784 694548 577020 694784
rect 577256 694548 577492 694784
rect 572560 694312 577492 694548
rect 572560 694076 572772 694312
rect 573008 694076 573244 694312
rect 573480 694076 573716 694312
rect 573952 694076 574188 694312
rect 574424 694076 574660 694312
rect 574896 694076 575132 694312
rect 575368 694076 575604 694312
rect 575840 694076 576076 694312
rect 576312 694076 576548 694312
rect 576784 694076 577020 694312
rect 577256 694076 577492 694312
rect 572560 693840 577492 694076
rect 572560 693604 572772 693840
rect 573008 693604 573244 693840
rect 573480 693604 573716 693840
rect 573952 693604 574188 693840
rect 574424 693604 574660 693840
rect 574896 693604 575132 693840
rect 575368 693604 575604 693840
rect 575840 693604 576076 693840
rect 576312 693604 576548 693840
rect 576784 693604 577020 693840
rect 577256 693604 577492 693840
rect 572560 693368 577492 693604
rect 572560 693132 572772 693368
rect 573008 693132 573244 693368
rect 573480 693132 573716 693368
rect 573952 693132 574188 693368
rect 574424 693132 574660 693368
rect 574896 693132 575132 693368
rect 575368 693132 575604 693368
rect 575840 693132 576076 693368
rect 576312 693132 576548 693368
rect 576784 693132 577020 693368
rect 577256 693132 577492 693368
rect 572560 692896 577492 693132
rect 572560 692660 572772 692896
rect 573008 692660 573244 692896
rect 573480 692660 573716 692896
rect 573952 692660 574188 692896
rect 574424 692660 574660 692896
rect 574896 692660 575132 692896
rect 575368 692660 575604 692896
rect 575840 692660 576076 692896
rect 576312 692660 576548 692896
rect 576784 692660 577020 692896
rect 577256 692660 577492 692896
rect 562456 644584 567424 654608
rect 562456 639784 562480 644584
rect 567400 639784 567424 644584
rect 562456 634584 567424 639784
rect 562456 629784 562480 634584
rect 567400 629784 567424 634584
rect 562456 522504 567424 629784
rect 562456 522268 562624 522504
rect 562860 522268 563096 522504
rect 563332 522268 563568 522504
rect 563804 522268 564040 522504
rect 564276 522268 564512 522504
rect 564748 522268 564984 522504
rect 565220 522268 565456 522504
rect 565692 522268 565928 522504
rect 566164 522268 566400 522504
rect 566636 522268 566872 522504
rect 567108 522268 567424 522504
rect 562456 522032 567424 522268
rect 562456 521796 562624 522032
rect 562860 521796 563096 522032
rect 563332 521796 563568 522032
rect 563804 521796 564040 522032
rect 564276 521796 564512 522032
rect 564748 521796 564984 522032
rect 565220 521796 565456 522032
rect 565692 521796 565928 522032
rect 566164 521796 566400 522032
rect 566636 521796 566872 522032
rect 567108 521796 567424 522032
rect 562456 521560 567424 521796
rect 562456 521324 562624 521560
rect 562860 521324 563096 521560
rect 563332 521324 563568 521560
rect 563804 521324 564040 521560
rect 564276 521324 564512 521560
rect 564748 521324 564984 521560
rect 565220 521324 565456 521560
rect 565692 521324 565928 521560
rect 566164 521324 566400 521560
rect 566636 521324 566872 521560
rect 567108 521324 567424 521560
rect 562456 521088 567424 521324
rect 562456 520852 562624 521088
rect 562860 520852 563096 521088
rect 563332 520852 563568 521088
rect 563804 520852 564040 521088
rect 564276 520852 564512 521088
rect 564748 520852 564984 521088
rect 565220 520852 565456 521088
rect 565692 520852 565928 521088
rect 566164 520852 566400 521088
rect 566636 520852 566872 521088
rect 567108 520852 567424 521088
rect 562456 520616 567424 520852
rect 562456 520380 562624 520616
rect 562860 520380 563096 520616
rect 563332 520380 563568 520616
rect 563804 520380 564040 520616
rect 564276 520380 564512 520616
rect 564748 520380 564984 520616
rect 565220 520380 565456 520616
rect 565692 520380 565928 520616
rect 566164 520380 566400 520616
rect 566636 520380 566872 520616
rect 567108 520380 567424 520616
rect 562456 520144 567424 520380
rect 562456 519908 562624 520144
rect 562860 519908 563096 520144
rect 563332 519908 563568 520144
rect 563804 519908 564040 520144
rect 564276 519908 564512 520144
rect 564748 519908 564984 520144
rect 565220 519908 565456 520144
rect 565692 519908 565928 520144
rect 566164 519908 566400 520144
rect 566636 519908 566872 520144
rect 567108 519908 567424 520144
rect 562456 519672 567424 519908
rect 562456 519436 562624 519672
rect 562860 519436 563096 519672
rect 563332 519436 563568 519672
rect 563804 519436 564040 519672
rect 564276 519436 564512 519672
rect 564748 519436 564984 519672
rect 565220 519436 565456 519672
rect 565692 519436 565928 519672
rect 566164 519436 566400 519672
rect 566636 519436 566872 519672
rect 567108 519436 567424 519672
rect 562456 519200 567424 519436
rect 562456 518964 562624 519200
rect 562860 518964 563096 519200
rect 563332 518964 563568 519200
rect 563804 518964 564040 519200
rect 564276 518964 564512 519200
rect 564748 518964 564984 519200
rect 565220 518964 565456 519200
rect 565692 518964 565928 519200
rect 566164 518964 566400 519200
rect 566636 518964 566872 519200
rect 567108 518964 567424 519200
rect 562456 518728 567424 518964
rect 562456 518492 562624 518728
rect 562860 518492 563096 518728
rect 563332 518492 563568 518728
rect 563804 518492 564040 518728
rect 564276 518492 564512 518728
rect 564748 518492 564984 518728
rect 565220 518492 565456 518728
rect 565692 518492 565928 518728
rect 566164 518492 566400 518728
rect 566636 518492 566872 518728
rect 567108 518492 567424 518728
rect 562456 518256 567424 518492
rect 562456 518020 562624 518256
rect 562860 518020 563096 518256
rect 563332 518020 563568 518256
rect 563804 518020 564040 518256
rect 564276 518020 564512 518256
rect 564748 518020 564984 518256
rect 565220 518020 565456 518256
rect 565692 518020 565928 518256
rect 566164 518020 566400 518256
rect 566636 518020 566872 518256
rect 567108 518020 567424 518256
rect 562456 517784 567424 518020
rect 562456 517548 562624 517784
rect 562860 517548 563096 517784
rect 563332 517548 563568 517784
rect 563804 517548 564040 517784
rect 564276 517548 564512 517784
rect 564748 517548 564984 517784
rect 565220 517548 565456 517784
rect 565692 517548 565928 517784
rect 566164 517548 566400 517784
rect 566636 517548 566872 517784
rect 567108 517548 567424 517784
rect 562456 517312 567424 517548
rect 562456 517076 562624 517312
rect 562860 517076 563096 517312
rect 563332 517076 563568 517312
rect 563804 517076 564040 517312
rect 564276 517076 564512 517312
rect 564748 517076 564984 517312
rect 565220 517076 565456 517312
rect 565692 517076 565928 517312
rect 566164 517076 566400 517312
rect 566636 517076 566872 517312
rect 567108 517076 567424 517312
rect 562456 516840 567424 517076
rect 562456 516604 562624 516840
rect 562860 516604 563096 516840
rect 563332 516604 563568 516840
rect 563804 516604 564040 516840
rect 564276 516604 564512 516840
rect 564748 516604 564984 516840
rect 565220 516604 565456 516840
rect 565692 516604 565928 516840
rect 566164 516604 566400 516840
rect 566636 516604 566872 516840
rect 567108 516604 567424 516840
rect 562456 495782 567424 516604
rect 562456 495546 562624 495782
rect 562860 495546 563096 495782
rect 563332 495546 563568 495782
rect 563804 495546 564040 495782
rect 564276 495546 564512 495782
rect 564748 495546 564984 495782
rect 565220 495546 565456 495782
rect 565692 495546 565928 495782
rect 566164 495546 566400 495782
rect 566636 495546 566872 495782
rect 567108 495546 567424 495782
rect 512174 472390 525651 472484
rect 512174 472070 518572 472390
rect 518892 472070 519272 472390
rect 519592 472070 519972 472390
rect 520292 472070 520672 472390
rect 520992 472070 521372 472390
rect 521692 472070 522072 472390
rect 522392 472070 522772 472390
rect 523092 472070 523472 472390
rect 523792 472070 524172 472390
rect 524492 472070 524872 472390
rect 525192 472070 525651 472390
rect 512174 471268 525651 472070
rect 512174 470948 518572 471268
rect 518892 470948 519272 471268
rect 519592 470948 519972 471268
rect 520292 470948 520672 471268
rect 520992 470948 521372 471268
rect 521692 470948 522072 471268
rect 522392 470948 522772 471268
rect 523092 470948 523472 471268
rect 523792 470948 524172 471268
rect 524492 470948 524872 471268
rect 525192 470948 525651 471268
rect 512174 470146 525651 470948
rect 512174 469826 518572 470146
rect 518892 469826 519272 470146
rect 519592 469826 519972 470146
rect 520292 469826 520672 470146
rect 520992 469826 521372 470146
rect 521692 469826 522072 470146
rect 522392 469826 522772 470146
rect 523092 469826 523472 470146
rect 523792 469826 524172 470146
rect 524492 469826 524872 470146
rect 525192 469826 525651 470146
rect 512174 469024 525651 469826
rect 512174 468704 518572 469024
rect 518892 468704 519272 469024
rect 519592 468704 519972 469024
rect 520292 468704 520672 469024
rect 520992 468704 521372 469024
rect 521692 468704 522072 469024
rect 522392 468704 522772 469024
rect 523092 468704 523472 469024
rect 523792 468704 524172 469024
rect 524492 468704 524872 469024
rect 525192 468704 525651 469024
rect 512174 467902 525651 468704
rect 512174 467582 518572 467902
rect 518892 467582 519272 467902
rect 519592 467582 519972 467902
rect 520292 467582 520672 467902
rect 520992 467582 521372 467902
rect 521692 467582 522072 467902
rect 522392 467582 522772 467902
rect 523092 467582 523472 467902
rect 523792 467582 524172 467902
rect 524492 467582 524872 467902
rect 525192 467582 525651 467902
rect 512174 466780 525651 467582
rect 512174 466460 518572 466780
rect 518892 466460 519272 466780
rect 519592 466460 519972 466780
rect 520292 466460 520672 466780
rect 520992 466460 521372 466780
rect 521692 466460 522072 466780
rect 522392 466460 522772 466780
rect 523092 466460 523472 466780
rect 523792 466460 524172 466780
rect 524492 466460 524872 466780
rect 525192 466460 525651 466780
rect 512174 465658 525651 466460
rect 512174 465338 518572 465658
rect 518892 465338 519272 465658
rect 519592 465338 519972 465658
rect 520292 465338 520672 465658
rect 520992 465338 521372 465658
rect 521692 465338 522072 465658
rect 522392 465338 522772 465658
rect 523092 465338 523472 465658
rect 523792 465338 524172 465658
rect 524492 465338 524872 465658
rect 525192 465338 525651 465658
rect 512174 464536 525651 465338
rect 512174 464216 518572 464536
rect 518892 464216 519272 464536
rect 519592 464216 519972 464536
rect 520292 464216 520672 464536
rect 520992 464216 521372 464536
rect 521692 464216 522072 464536
rect 522392 464216 522772 464536
rect 523092 464216 523472 464536
rect 523792 464216 524172 464536
rect 524492 464216 524872 464536
rect 525192 464216 525651 464536
rect 512174 463414 525651 464216
rect 512174 463094 518572 463414
rect 518892 463094 519272 463414
rect 519592 463094 519972 463414
rect 520292 463094 520672 463414
rect 520992 463094 521372 463414
rect 521692 463094 522072 463414
rect 522392 463094 522772 463414
rect 523092 463094 523472 463414
rect 523792 463094 524172 463414
rect 524492 463094 524872 463414
rect 525192 463094 525651 463414
rect 512174 462292 525651 463094
rect 512174 461972 518572 462292
rect 518892 461972 519272 462292
rect 519592 461972 519972 462292
rect 520292 461972 520672 462292
rect 520992 461972 521372 462292
rect 521692 461972 522072 462292
rect 522392 461972 522772 462292
rect 523092 461972 523472 462292
rect 523792 461972 524172 462292
rect 524492 461972 524872 462292
rect 525192 461972 525651 462292
rect 512174 460198 525651 461972
rect 512136 439888 512234 460198
rect 513206 439888 525651 460198
rect 512136 439870 525651 439888
rect 562456 455480 567424 495546
rect 562456 455244 562624 455480
rect 562860 455244 563096 455480
rect 563332 455244 563568 455480
rect 563804 455244 564040 455480
rect 564276 455244 564512 455480
rect 564748 455244 564984 455480
rect 565220 455244 565456 455480
rect 565692 455244 565928 455480
rect 566164 455244 566400 455480
rect 566636 455244 566872 455480
rect 567108 455244 567424 455480
rect 512136 439714 525376 439870
rect 562456 377364 567424 455244
rect 562456 377128 562624 377364
rect 562860 377128 563096 377364
rect 563332 377128 563568 377364
rect 563804 377128 564040 377364
rect 564276 377128 564512 377364
rect 564748 377128 564984 377364
rect 565220 377128 565456 377364
rect 565692 377128 565928 377364
rect 566164 377128 566400 377364
rect 566636 377128 566872 377364
rect 567108 377128 567424 377364
rect 562456 376892 567424 377128
rect 562456 376656 562624 376892
rect 562860 376656 563096 376892
rect 563332 376656 563568 376892
rect 563804 376656 564040 376892
rect 564276 376656 564512 376892
rect 564748 376656 564984 376892
rect 565220 376656 565456 376892
rect 565692 376656 565928 376892
rect 566164 376656 566400 376892
rect 566636 376656 566872 376892
rect 567108 376656 567424 376892
rect 562456 376420 567424 376656
rect 562456 376184 562624 376420
rect 562860 376184 563096 376420
rect 563332 376184 563568 376420
rect 563804 376184 564040 376420
rect 564276 376184 564512 376420
rect 564748 376184 564984 376420
rect 565220 376184 565456 376420
rect 565692 376184 565928 376420
rect 566164 376184 566400 376420
rect 566636 376184 566872 376420
rect 567108 376184 567424 376420
rect 562456 375948 567424 376184
rect 562456 375712 562624 375948
rect 562860 375712 563096 375948
rect 563332 375712 563568 375948
rect 563804 375712 564040 375948
rect 564276 375712 564512 375948
rect 564748 375712 564984 375948
rect 565220 375712 565456 375948
rect 565692 375712 565928 375948
rect 566164 375712 566400 375948
rect 566636 375712 566872 375948
rect 567108 375712 567424 375948
rect 562456 375476 567424 375712
rect 562456 375240 562624 375476
rect 562860 375240 563096 375476
rect 563332 375240 563568 375476
rect 563804 375240 564040 375476
rect 564276 375240 564512 375476
rect 564748 375240 564984 375476
rect 565220 375240 565456 375476
rect 565692 375240 565928 375476
rect 566164 375240 566400 375476
rect 566636 375240 566872 375476
rect 567108 375240 567424 375476
rect 562456 375004 567424 375240
rect 562456 374768 562624 375004
rect 562860 374768 563096 375004
rect 563332 374768 563568 375004
rect 563804 374768 564040 375004
rect 564276 374768 564512 375004
rect 564748 374768 564984 375004
rect 565220 374768 565456 375004
rect 565692 374768 565928 375004
rect 566164 374768 566400 375004
rect 566636 374768 566872 375004
rect 567108 374768 567424 375004
rect 562456 374532 567424 374768
rect 562456 374296 562624 374532
rect 562860 374296 563096 374532
rect 563332 374296 563568 374532
rect 563804 374296 564040 374532
rect 564276 374296 564512 374532
rect 564748 374296 564984 374532
rect 565220 374296 565456 374532
rect 565692 374296 565928 374532
rect 566164 374296 566400 374532
rect 566636 374296 566872 374532
rect 567108 374296 567424 374532
rect 562456 374060 567424 374296
rect 562456 373824 562624 374060
rect 562860 373824 563096 374060
rect 563332 373824 563568 374060
rect 563804 373824 564040 374060
rect 564276 373824 564512 374060
rect 564748 373824 564984 374060
rect 565220 373824 565456 374060
rect 565692 373824 565928 374060
rect 566164 373824 566400 374060
rect 566636 373824 566872 374060
rect 567108 373824 567424 374060
rect 562456 373588 567424 373824
rect 562456 373352 562624 373588
rect 562860 373352 563096 373588
rect 563332 373352 563568 373588
rect 563804 373352 564040 373588
rect 564276 373352 564512 373588
rect 564748 373352 564984 373588
rect 565220 373352 565456 373588
rect 565692 373352 565928 373588
rect 566164 373352 566400 373588
rect 566636 373352 566872 373588
rect 567108 373352 567424 373588
rect 562456 373116 567424 373352
rect 562456 372880 562624 373116
rect 562860 372880 563096 373116
rect 563332 372880 563568 373116
rect 563804 372880 564040 373116
rect 564276 372880 564512 373116
rect 564748 372880 564984 373116
rect 565220 372880 565456 373116
rect 565692 372880 565928 373116
rect 566164 372880 566400 373116
rect 566636 372880 566872 373116
rect 567108 372880 567424 373116
rect 562456 372644 567424 372880
rect 562456 372408 562624 372644
rect 562860 372408 563096 372644
rect 563332 372408 563568 372644
rect 563804 372408 564040 372644
rect 564276 372408 564512 372644
rect 564748 372408 564984 372644
rect 565220 372408 565456 372644
rect 565692 372408 565928 372644
rect 566164 372408 566400 372644
rect 566636 372408 566872 372644
rect 567108 372408 567424 372644
rect 562456 372172 567424 372408
rect 562456 371936 562624 372172
rect 562860 371936 563096 372172
rect 563332 371936 563568 372172
rect 563804 371936 564040 372172
rect 564276 371936 564512 372172
rect 564748 371936 564984 372172
rect 565220 371936 565456 372172
rect 565692 371936 565928 372172
rect 566164 371936 566400 372172
rect 566636 371936 566872 372172
rect 567108 371936 567424 372172
rect 562456 371700 567424 371936
rect 562456 371464 562624 371700
rect 562860 371464 563096 371700
rect 563332 371464 563568 371700
rect 563804 371464 564040 371700
rect 564276 371464 564512 371700
rect 564748 371464 564984 371700
rect 565220 371464 565456 371700
rect 565692 371464 565928 371700
rect 566164 371464 566400 371700
rect 566636 371464 566872 371700
rect 567108 371464 567424 371700
rect 562456 303322 567424 371464
rect 572560 495782 577480 692660
rect 572560 495546 572784 495782
rect 573020 495546 573256 495782
rect 573492 495546 573728 495782
rect 573964 495546 574200 495782
rect 574436 495546 574672 495782
rect 574908 495546 575144 495782
rect 575380 495546 575616 495782
rect 575852 495546 576088 495782
rect 576324 495546 576560 495782
rect 576796 495546 577032 495782
rect 577268 495546 577480 495782
rect 572560 484272 577480 495546
rect 572560 484036 577492 484272
rect 572560 483800 572772 484036
rect 573008 483800 573244 484036
rect 573480 483800 573716 484036
rect 573952 483800 574188 484036
rect 574424 483800 574660 484036
rect 574896 483800 575132 484036
rect 575368 483800 575604 484036
rect 575840 483800 576076 484036
rect 576312 483800 576548 484036
rect 576784 483800 577020 484036
rect 577256 483800 577492 484036
rect 572560 483564 577492 483800
rect 572560 483328 572772 483564
rect 573008 483328 573244 483564
rect 573480 483328 573716 483564
rect 573952 483328 574188 483564
rect 574424 483328 574660 483564
rect 574896 483328 575132 483564
rect 575368 483328 575604 483564
rect 575840 483328 576076 483564
rect 576312 483328 576548 483564
rect 576784 483328 577020 483564
rect 577256 483328 577492 483564
rect 572560 483092 577492 483328
rect 572560 482856 572772 483092
rect 573008 482856 573244 483092
rect 573480 482856 573716 483092
rect 573952 482856 574188 483092
rect 574424 482856 574660 483092
rect 574896 482856 575132 483092
rect 575368 482856 575604 483092
rect 575840 482856 576076 483092
rect 576312 482856 576548 483092
rect 576784 482856 577020 483092
rect 577256 482856 577492 483092
rect 572560 482620 577492 482856
rect 572560 482384 572772 482620
rect 573008 482384 573244 482620
rect 573480 482384 573716 482620
rect 573952 482384 574188 482620
rect 574424 482384 574660 482620
rect 574896 482384 575132 482620
rect 575368 482384 575604 482620
rect 575840 482384 576076 482620
rect 576312 482384 576548 482620
rect 576784 482384 577020 482620
rect 577256 482384 577492 482620
rect 572560 482148 577492 482384
rect 572560 481912 572772 482148
rect 573008 481912 573244 482148
rect 573480 481912 573716 482148
rect 573952 481912 574188 482148
rect 574424 481912 574660 482148
rect 574896 481912 575132 482148
rect 575368 481912 575604 482148
rect 575840 481912 576076 482148
rect 576312 481912 576548 482148
rect 576784 481912 577020 482148
rect 577256 481912 577492 482148
rect 572560 481676 577492 481912
rect 572560 481440 572772 481676
rect 573008 481440 573244 481676
rect 573480 481440 573716 481676
rect 573952 481440 574188 481676
rect 574424 481440 574660 481676
rect 574896 481440 575132 481676
rect 575368 481440 575604 481676
rect 575840 481440 576076 481676
rect 576312 481440 576548 481676
rect 576784 481440 577020 481676
rect 577256 481440 577492 481676
rect 572560 481204 577492 481440
rect 572560 480968 572772 481204
rect 573008 480968 573244 481204
rect 573480 480968 573716 481204
rect 573952 480968 574188 481204
rect 574424 480968 574660 481204
rect 574896 480968 575132 481204
rect 575368 480968 575604 481204
rect 575840 480968 576076 481204
rect 576312 480968 576548 481204
rect 576784 480968 577020 481204
rect 577256 480968 577492 481204
rect 572560 480732 577492 480968
rect 572560 480496 572772 480732
rect 573008 480496 573244 480732
rect 573480 480496 573716 480732
rect 573952 480496 574188 480732
rect 574424 480496 574660 480732
rect 574896 480496 575132 480732
rect 575368 480496 575604 480732
rect 575840 480496 576076 480732
rect 576312 480496 576548 480732
rect 576784 480496 577020 480732
rect 577256 480496 577492 480732
rect 572560 480260 577492 480496
rect 572560 480024 572772 480260
rect 573008 480024 573244 480260
rect 573480 480024 573716 480260
rect 573952 480024 574188 480260
rect 574424 480024 574660 480260
rect 574896 480024 575132 480260
rect 575368 480024 575604 480260
rect 575840 480024 576076 480260
rect 576312 480024 576548 480260
rect 576784 480024 577020 480260
rect 577256 480024 577492 480260
rect 572560 479788 577492 480024
rect 572560 479552 572772 479788
rect 573008 479552 573244 479788
rect 573480 479552 573716 479788
rect 573952 479552 574188 479788
rect 574424 479552 574660 479788
rect 574896 479552 575132 479788
rect 575368 479552 575604 479788
rect 575840 479552 576076 479788
rect 576312 479552 576548 479788
rect 576784 479552 577020 479788
rect 577256 479552 577492 479788
rect 572560 479316 577492 479552
rect 572560 479080 572772 479316
rect 573008 479080 573244 479316
rect 573480 479080 573716 479316
rect 573952 479080 574188 479316
rect 574424 479080 574660 479316
rect 574896 479080 575132 479316
rect 575368 479080 575604 479316
rect 575840 479080 576076 479316
rect 576312 479080 576548 479316
rect 576784 479080 577020 479316
rect 577256 479080 577492 479316
rect 572560 478844 577492 479080
rect 572560 478608 572772 478844
rect 573008 478608 573244 478844
rect 573480 478608 573716 478844
rect 573952 478608 574188 478844
rect 574424 478608 574660 478844
rect 574896 478608 575132 478844
rect 575368 478608 575604 478844
rect 575840 478608 576076 478844
rect 576312 478608 576548 478844
rect 576784 478608 577020 478844
rect 577256 478608 577492 478844
rect 572560 478372 577492 478608
rect 572560 478136 572772 478372
rect 573008 478136 573244 478372
rect 573480 478136 573716 478372
rect 573952 478136 574188 478372
rect 574424 478136 574660 478372
rect 574896 478136 575132 478372
rect 575368 478136 575604 478372
rect 575840 478136 576076 478372
rect 576312 478136 576548 478372
rect 576784 478136 577020 478372
rect 577256 478136 577492 478372
rect 572560 477900 577492 478136
rect 572560 477664 572772 477900
rect 573008 477664 573244 477900
rect 573480 477664 573716 477900
rect 573952 477664 574188 477900
rect 574424 477664 574660 477900
rect 574896 477664 575132 477900
rect 575368 477664 575604 477900
rect 575840 477664 576076 477900
rect 576312 477664 576548 477900
rect 576784 477664 577020 477900
rect 577256 477664 577492 477900
rect 572560 455480 577480 477664
rect 572560 455244 572784 455480
rect 573020 455244 573256 455480
rect 573492 455244 573728 455480
rect 573964 455244 574200 455480
rect 574436 455244 574672 455480
rect 574908 455244 575144 455480
rect 575380 455244 575616 455480
rect 575852 455244 576088 455480
rect 576324 455244 576560 455480
rect 576796 455244 577032 455480
rect 577268 455244 577480 455480
rect 572560 426924 577480 455244
rect 572560 426688 577492 426924
rect 572560 426452 572772 426688
rect 573008 426452 573244 426688
rect 573480 426452 573716 426688
rect 573952 426452 574188 426688
rect 574424 426452 574660 426688
rect 574896 426452 575132 426688
rect 575368 426452 575604 426688
rect 575840 426452 576076 426688
rect 576312 426452 576548 426688
rect 576784 426452 577020 426688
rect 577256 426452 577492 426688
rect 572560 426216 577492 426452
rect 572560 425980 572772 426216
rect 573008 425980 573244 426216
rect 573480 425980 573716 426216
rect 573952 425980 574188 426216
rect 574424 425980 574660 426216
rect 574896 425980 575132 426216
rect 575368 425980 575604 426216
rect 575840 425980 576076 426216
rect 576312 425980 576548 426216
rect 576784 425980 577020 426216
rect 577256 425980 577492 426216
rect 572560 425744 577492 425980
rect 572560 425508 572772 425744
rect 573008 425508 573244 425744
rect 573480 425508 573716 425744
rect 573952 425508 574188 425744
rect 574424 425508 574660 425744
rect 574896 425508 575132 425744
rect 575368 425508 575604 425744
rect 575840 425508 576076 425744
rect 576312 425508 576548 425744
rect 576784 425508 577020 425744
rect 577256 425508 577492 425744
rect 572560 425272 577492 425508
rect 572560 425036 572772 425272
rect 573008 425036 573244 425272
rect 573480 425036 573716 425272
rect 573952 425036 574188 425272
rect 574424 425036 574660 425272
rect 574896 425036 575132 425272
rect 575368 425036 575604 425272
rect 575840 425036 576076 425272
rect 576312 425036 576548 425272
rect 576784 425036 577020 425272
rect 577256 425036 577492 425272
rect 572560 424800 577492 425036
rect 572560 424564 572772 424800
rect 573008 424564 573244 424800
rect 573480 424564 573716 424800
rect 573952 424564 574188 424800
rect 574424 424564 574660 424800
rect 574896 424564 575132 424800
rect 575368 424564 575604 424800
rect 575840 424564 576076 424800
rect 576312 424564 576548 424800
rect 576784 424564 577020 424800
rect 577256 424564 577492 424800
rect 572560 424328 577492 424564
rect 572560 424092 572772 424328
rect 573008 424092 573244 424328
rect 573480 424092 573716 424328
rect 573952 424092 574188 424328
rect 574424 424092 574660 424328
rect 574896 424092 575132 424328
rect 575368 424092 575604 424328
rect 575840 424092 576076 424328
rect 576312 424092 576548 424328
rect 576784 424092 577020 424328
rect 577256 424092 577492 424328
rect 572560 423856 577492 424092
rect 572560 423620 572772 423856
rect 573008 423620 573244 423856
rect 573480 423620 573716 423856
rect 573952 423620 574188 423856
rect 574424 423620 574660 423856
rect 574896 423620 575132 423856
rect 575368 423620 575604 423856
rect 575840 423620 576076 423856
rect 576312 423620 576548 423856
rect 576784 423620 577020 423856
rect 577256 423620 577492 423856
rect 572560 423384 577492 423620
rect 572560 423148 572772 423384
rect 573008 423148 573244 423384
rect 573480 423148 573716 423384
rect 573952 423148 574188 423384
rect 574424 423148 574660 423384
rect 574896 423148 575132 423384
rect 575368 423148 575604 423384
rect 575840 423148 576076 423384
rect 576312 423148 576548 423384
rect 576784 423148 577020 423384
rect 577256 423148 577492 423384
rect 572560 422912 577492 423148
rect 572560 422676 572772 422912
rect 573008 422676 573244 422912
rect 573480 422676 573716 422912
rect 573952 422676 574188 422912
rect 574424 422676 574660 422912
rect 574896 422676 575132 422912
rect 575368 422676 575604 422912
rect 575840 422676 576076 422912
rect 576312 422676 576548 422912
rect 576784 422676 577020 422912
rect 577256 422676 577492 422912
rect 572560 422440 577492 422676
rect 572560 422204 572772 422440
rect 573008 422204 573244 422440
rect 573480 422204 573716 422440
rect 573952 422204 574188 422440
rect 574424 422204 574660 422440
rect 574896 422204 575132 422440
rect 575368 422204 575604 422440
rect 575840 422204 576076 422440
rect 576312 422204 576548 422440
rect 576784 422204 577020 422440
rect 577256 422204 577492 422440
rect 572560 421968 577492 422204
rect 572560 421732 572772 421968
rect 573008 421732 573244 421968
rect 573480 421732 573716 421968
rect 573952 421732 574188 421968
rect 574424 421732 574660 421968
rect 574896 421732 575132 421968
rect 575368 421732 575604 421968
rect 575840 421732 576076 421968
rect 576312 421732 576548 421968
rect 576784 421732 577020 421968
rect 577256 421732 577492 421968
rect 572560 421496 577492 421732
rect 572560 421260 572772 421496
rect 573008 421260 573244 421496
rect 573480 421260 573716 421496
rect 573952 421260 574188 421496
rect 574424 421260 574660 421496
rect 574896 421260 575132 421496
rect 575368 421260 575604 421496
rect 575840 421260 576076 421496
rect 576312 421260 576548 421496
rect 576784 421260 577020 421496
rect 577256 421260 577492 421496
rect 572560 421024 577492 421260
rect 572560 420788 572772 421024
rect 573008 420788 573244 421024
rect 573480 420788 573716 421024
rect 573952 420788 574188 421024
rect 574424 420788 574660 421024
rect 574896 420788 575132 421024
rect 575368 420788 575604 421024
rect 575840 420788 576076 421024
rect 576312 420788 576548 421024
rect 576784 420788 577020 421024
rect 577256 420788 577492 421024
rect 572560 420552 577492 420788
rect 572560 420316 572772 420552
rect 573008 420316 573244 420552
rect 573480 420316 573716 420552
rect 573952 420316 574188 420552
rect 574424 420316 574660 420552
rect 574896 420316 575132 420552
rect 575368 420316 575604 420552
rect 575840 420316 576076 420552
rect 576312 420316 576548 420552
rect 576784 420316 577020 420552
rect 577256 420316 577492 420552
rect 572560 312500 577480 420316
<< comment >>
rect -100 704000 584100 704100
rect -100 0 0 704000
rect 584000 0 584100 704000
rect -100 -100 584100 0
<< res2p85 >>
rect 518276 459312 521604 459886
rect 518276 458494 521604 459068
rect 518276 457676 521604 458250
rect 518686 456040 522990 456614
rect 518686 455222 522990 455796
rect 518686 454404 522990 454978
rect 518686 453586 522990 454160
rect 516620 451132 522928 451706
rect 516620 450314 522928 450888
rect 516620 449496 522928 450070
rect 516620 448678 522928 449252
rect 516620 447860 522928 448434
rect 516620 447042 522928 447616
rect 516620 446224 522928 446798
rect 516620 445406 522928 445980
rect 516620 444588 522928 445162
rect 516620 443770 522928 444344
rect 516620 442952 522928 443526
rect 516620 442134 522928 442708
rect 516620 441316 522928 441890
rect 516620 440498 522928 441072
rect 516620 439680 522928 440254
rect 516620 438862 522928 439436
rect 516620 438044 522928 438618
<< pnp3p40 >>
rect 503497 437321 504531 438355
rect 504785 437321 505819 438355
rect 506073 437321 507107 438355
rect 507361 437321 508395 438355
rect 508649 437321 509683 438355
rect 509937 437321 510971 438355
rect 511225 437321 512259 438355
rect 512513 437321 513547 438355
rect 503497 436033 504531 437067
rect 504785 436033 505819 437067
rect 506073 436033 507107 437067
rect 507361 436033 508395 437067
rect 508649 436033 509683 437067
rect 509937 436033 510971 437067
rect 511225 436033 512259 437067
rect 512513 436033 513547 437067
rect 503497 434745 504531 435779
rect 504785 434745 505819 435779
rect 506073 434745 507107 435779
rect 507361 434745 508395 435779
rect 508649 434745 509683 435779
rect 509937 434745 510971 435779
rect 511225 434745 512259 435779
rect 512513 434745 513547 435779
rect 503497 433457 504531 434491
rect 504785 433457 505819 434491
rect 506073 433457 507107 434491
rect 507361 433457 508395 434491
rect 508649 433457 509683 434491
rect 509937 433457 510971 434491
rect 511225 433457 512259 434491
rect 512513 433457 513547 434491
rect 503497 432169 504531 433203
rect 504785 432169 505819 433203
rect 506073 432169 507107 433203
rect 507361 432169 508395 433203
rect 508649 432169 509683 433203
rect 509937 432169 510971 433203
rect 511225 432169 512259 433203
rect 512513 432169 513547 433203
<< labels >>
flabel metal3 s 583520 269230 584800 269342 0 FreeSans 1120 0 0 0 gpio_analog[0]
port 0 nsew signal bidirectional
flabel metal3 s -800 381864 480 381976 0 FreeSans 1120 0 0 0 gpio_analog[10]
port 1 nsew signal bidirectional
flabel metal3 s -800 338642 480 338754 0 FreeSans 1120 0 0 0 gpio_analog[11]
port 2 nsew signal bidirectional
flabel metal3 s -800 295420 480 295532 0 FreeSans 1120 0 0 0 gpio_analog[12]
port 3 nsew signal bidirectional
flabel metal3 s -800 252398 480 252510 0 FreeSans 1120 0 0 0 gpio_analog[13]
port 4 nsew signal bidirectional
flabel metal3 s -800 124776 480 124888 0 FreeSans 1120 0 0 0 gpio_analog[14]
port 5 nsew signal bidirectional
flabel metal3 s -800 81554 480 81666 0 FreeSans 1120 0 0 0 gpio_analog[15]
port 6 nsew signal bidirectional
flabel metal3 s -800 38332 480 38444 0 FreeSans 1120 0 0 0 gpio_analog[16]
port 7 nsew signal bidirectional
flabel metal3 s -800 16910 480 17022 0 FreeSans 1120 0 0 0 gpio_analog[17]
port 8 nsew signal bidirectional
flabel metal3 s 583520 313652 584800 313764 0 FreeSans 1120 0 0 0 gpio_analog[1]
port 9 nsew signal bidirectional
flabel metal3 s 583520 358874 584800 358986 0 FreeSans 1120 0 0 0 gpio_analog[2]
port 10 nsew signal bidirectional
flabel metal3 s 583520 405296 584800 405408 0 FreeSans 1120 0 0 0 gpio_analog[3]
port 11 nsew signal bidirectional
flabel metal3 s 583520 449718 584800 449830 0 FreeSans 1120 0 0 0 gpio_analog[4]
port 12 nsew signal bidirectional
flabel metal3 s 583520 494140 584800 494252 0 FreeSans 1120 0 0 0 gpio_analog[5]
port 13 nsew signal bidirectional
flabel metal3 s 583520 583562 584800 583674 0 FreeSans 1120 0 0 0 gpio_analog[6]
port 14 nsew signal bidirectional
flabel metal3 s -800 511530 480 511642 0 FreeSans 1120 0 0 0 gpio_analog[7]
port 15 nsew signal bidirectional
flabel metal3 s -800 468308 480 468420 0 FreeSans 1120 0 0 0 gpio_analog[8]
port 16 nsew signal bidirectional
flabel metal3 s -800 425086 480 425198 0 FreeSans 1120 0 0 0 gpio_analog[9]
port 17 nsew signal bidirectional
flabel metal3 s 583520 270412 584800 270524 0 FreeSans 1120 0 0 0 gpio_noesd[0]
port 18 nsew signal bidirectional
flabel metal3 s -800 380682 480 380794 0 FreeSans 1120 0 0 0 gpio_noesd[10]
port 19 nsew signal bidirectional
flabel metal3 s -800 337460 480 337572 0 FreeSans 1120 0 0 0 gpio_noesd[11]
port 20 nsew signal bidirectional
flabel metal3 s -800 294238 480 294350 0 FreeSans 1120 0 0 0 gpio_noesd[12]
port 21 nsew signal bidirectional
flabel metal3 s -800 251216 480 251328 0 FreeSans 1120 0 0 0 gpio_noesd[13]
port 22 nsew signal bidirectional
flabel metal3 s -800 123594 480 123706 0 FreeSans 1120 0 0 0 gpio_noesd[14]
port 23 nsew signal bidirectional
flabel metal3 s -800 80372 480 80484 0 FreeSans 1120 0 0 0 gpio_noesd[15]
port 24 nsew signal bidirectional
flabel metal3 s -800 37150 480 37262 0 FreeSans 1120 0 0 0 gpio_noesd[16]
port 25 nsew signal bidirectional
flabel metal3 s -800 15728 480 15840 0 FreeSans 1120 0 0 0 gpio_noesd[17]
port 26 nsew signal bidirectional
flabel metal3 s 583520 314834 584800 314946 0 FreeSans 1120 0 0 0 gpio_noesd[1]
port 27 nsew signal bidirectional
flabel metal3 s 583520 360056 584800 360168 0 FreeSans 1120 0 0 0 gpio_noesd[2]
port 28 nsew signal bidirectional
flabel metal3 s 583520 406478 584800 406590 0 FreeSans 1120 0 0 0 gpio_noesd[3]
port 29 nsew signal bidirectional
flabel metal3 s 583520 450900 584800 451012 0 FreeSans 1120 0 0 0 gpio_noesd[4]
port 30 nsew signal bidirectional
flabel metal3 s 583520 495322 584800 495434 0 FreeSans 1120 0 0 0 gpio_noesd[5]
port 31 nsew signal bidirectional
flabel metal3 s 583520 584744 584800 584856 0 FreeSans 1120 0 0 0 gpio_noesd[6]
port 32 nsew signal bidirectional
flabel metal3 s -800 510348 480 510460 0 FreeSans 1120 0 0 0 gpio_noesd[7]
port 33 nsew signal bidirectional
flabel metal3 s -800 467126 480 467238 0 FreeSans 1120 0 0 0 gpio_noesd[8]
port 34 nsew signal bidirectional
flabel metal3 s -800 423904 480 424016 0 FreeSans 1120 0 0 0 gpio_noesd[9]
port 35 nsew signal bidirectional
flabel metal3 s 582300 677984 584800 682984 0 FreeSans 1120 0 0 0 io_analog[0]
port 36 nsew signal bidirectional
flabel metal3 s 0 680242 1700 685242 0 FreeSans 1120 0 0 0 io_analog[10]
port 37 nsew signal bidirectional
flabel metal3 s 566594 702300 571594 704800 0 FreeSans 1920 180 0 0 io_analog[1]
port 38 nsew signal bidirectional
flabel metal3 s 465394 702300 470394 704800 0 FreeSans 1920 180 0 0 io_analog[2]
port 39 nsew signal bidirectional
flabel metal3 s 413394 702300 418394 704800 0 FreeSans 1920 180 0 0 io_analog[3]
port 40 nsew signal bidirectional
flabel metal3 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal3 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal3 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal3 s 120194 702300 125194 704800 0 FreeSans 1920 180 0 0 io_analog[7]
port 44 nsew signal bidirectional
flabel metal3 s 68194 702300 73194 704800 0 FreeSans 1920 180 0 0 io_analog[8]
port 45 nsew signal bidirectional
flabel metal3 s 16194 702300 21194 704800 0 FreeSans 1920 180 0 0 io_analog[9]
port 46 nsew signal bidirectional
flabel metal3 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal3 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal3 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal3 s 326794 702300 328994 704800 0 FreeSans 1920 180 0 0 io_clamp_high[0]
port 50 nsew signal bidirectional
flabel metal3 s 225094 702300 227294 704800 0 FreeSans 1920 180 0 0 io_clamp_high[1]
port 51 nsew signal bidirectional
flabel metal3 s 173394 702300 175594 704800 0 FreeSans 1920 180 0 0 io_clamp_high[2]
port 52 nsew signal bidirectional
flabel metal3 s 324294 702300 326494 704800 0 FreeSans 1920 180 0 0 io_clamp_low[0]
port 53 nsew signal bidirectional
flabel metal3 s 222594 702300 224794 704800 0 FreeSans 1920 180 0 0 io_clamp_low[1]
port 54 nsew signal bidirectional
flabel metal3 s 170894 702300 173094 704800 0 FreeSans 1920 180 0 0 io_clamp_low[2]
port 55 nsew signal bidirectional
flabel metal3 s 583520 2726 584800 2838 0 FreeSans 1120 0 0 0 io_in[0]
port 56 nsew signal input
flabel metal3 s 583520 408842 584800 408954 0 FreeSans 1120 0 0 0 io_in[10]
port 57 nsew signal input
flabel metal3 s 583520 453264 584800 453376 0 FreeSans 1120 0 0 0 io_in[11]
port 58 nsew signal input
flabel metal3 s 583520 497686 584800 497798 0 FreeSans 1120 0 0 0 io_in[12]
port 59 nsew signal input
flabel metal3 s 583520 587108 584800 587220 0 FreeSans 1120 0 0 0 io_in[13]
port 60 nsew signal input
flabel metal3 s -800 507984 480 508096 0 FreeSans 1120 0 0 0 io_in[14]
port 61 nsew signal input
flabel metal3 s -800 464762 480 464874 0 FreeSans 1120 0 0 0 io_in[15]
port 62 nsew signal input
flabel metal3 s -800 421540 480 421652 0 FreeSans 1120 0 0 0 io_in[16]
port 63 nsew signal input
flabel metal3 s -800 378318 480 378430 0 FreeSans 1120 0 0 0 io_in[17]
port 64 nsew signal input
flabel metal3 s -800 335096 480 335208 0 FreeSans 1120 0 0 0 io_in[18]
port 65 nsew signal input
flabel metal3 s -800 291874 480 291986 0 FreeSans 1120 0 0 0 io_in[19]
port 66 nsew signal input
flabel metal3 s 583520 7454 584800 7566 0 FreeSans 1120 0 0 0 io_in[1]
port 67 nsew signal input
flabel metal3 s -800 248852 480 248964 0 FreeSans 1120 0 0 0 io_in[20]
port 68 nsew signal input
flabel metal3 s -800 121230 480 121342 0 FreeSans 1120 0 0 0 io_in[21]
port 69 nsew signal input
flabel metal3 s -800 78008 480 78120 0 FreeSans 1120 0 0 0 io_in[22]
port 70 nsew signal input
flabel metal3 s -800 34786 480 34898 0 FreeSans 1120 0 0 0 io_in[23]
port 71 nsew signal input
flabel metal3 s -800 13364 480 13476 0 FreeSans 1120 0 0 0 io_in[24]
port 72 nsew signal input
flabel metal3 s -800 8636 480 8748 0 FreeSans 1120 0 0 0 io_in[25]
port 73 nsew signal input
flabel metal3 s -800 3908 480 4020 0 FreeSans 1120 0 0 0 io_in[26]
port 74 nsew signal input
flabel metal3 s 583520 12182 584800 12294 0 FreeSans 1120 0 0 0 io_in[2]
port 75 nsew signal input
flabel metal3 s 583520 16910 584800 17022 0 FreeSans 1120 0 0 0 io_in[3]
port 76 nsew signal input
flabel metal3 s 583520 21638 584800 21750 0 FreeSans 1120 0 0 0 io_in[4]
port 77 nsew signal input
flabel metal3 s 583520 48096 584800 48208 0 FreeSans 1120 0 0 0 io_in[5]
port 78 nsew signal input
flabel metal3 s 583520 92754 584800 92866 0 FreeSans 1120 0 0 0 io_in[6]
port 79 nsew signal input
flabel metal3 s 583520 272776 584800 272888 0 FreeSans 1120 0 0 0 io_in[7]
port 80 nsew signal input
flabel metal3 s 583520 317198 584800 317310 0 FreeSans 1120 0 0 0 io_in[8]
port 81 nsew signal input
flabel metal3 s 583520 362420 584800 362532 0 FreeSans 1120 0 0 0 io_in[9]
port 82 nsew signal input
flabel metal3 s 583520 1544 584800 1656 0 FreeSans 1120 0 0 0 io_in_3v3[0]
port 83 nsew signal input
flabel metal3 s 583520 407660 584800 407772 0 FreeSans 1120 0 0 0 io_in_3v3[10]
port 84 nsew signal input
flabel metal3 s 583520 452082 584800 452194 0 FreeSans 1120 0 0 0 io_in_3v3[11]
port 85 nsew signal input
flabel metal3 s 583520 496504 584800 496616 0 FreeSans 1120 0 0 0 io_in_3v3[12]
port 86 nsew signal input
flabel metal3 s 583520 585926 584800 586038 0 FreeSans 1120 0 0 0 io_in_3v3[13]
port 87 nsew signal input
flabel metal3 s -800 509166 480 509278 0 FreeSans 1120 0 0 0 io_in_3v3[14]
port 88 nsew signal input
flabel metal3 s -800 465944 480 466056 0 FreeSans 1120 0 0 0 io_in_3v3[15]
port 89 nsew signal input
flabel metal3 s -800 422722 480 422834 0 FreeSans 1120 0 0 0 io_in_3v3[16]
port 90 nsew signal input
flabel metal3 s -800 379500 480 379612 0 FreeSans 1120 0 0 0 io_in_3v3[17]
port 91 nsew signal input
flabel metal3 s -800 336278 480 336390 0 FreeSans 1120 0 0 0 io_in_3v3[18]
port 92 nsew signal input
flabel metal3 s -800 293056 480 293168 0 FreeSans 1120 0 0 0 io_in_3v3[19]
port 93 nsew signal input
flabel metal3 s 583520 6272 584800 6384 0 FreeSans 1120 0 0 0 io_in_3v3[1]
port 94 nsew signal input
flabel metal3 s -800 250034 480 250146 0 FreeSans 1120 0 0 0 io_in_3v3[20]
port 95 nsew signal input
flabel metal3 s -800 122412 480 122524 0 FreeSans 1120 0 0 0 io_in_3v3[21]
port 96 nsew signal input
flabel metal3 s -800 79190 480 79302 0 FreeSans 1120 0 0 0 io_in_3v3[22]
port 97 nsew signal input
flabel metal3 s -800 35968 480 36080 0 FreeSans 1120 0 0 0 io_in_3v3[23]
port 98 nsew signal input
flabel metal3 s -800 14546 480 14658 0 FreeSans 1120 0 0 0 io_in_3v3[24]
port 99 nsew signal input
flabel metal3 s -800 9818 480 9930 0 FreeSans 1120 0 0 0 io_in_3v3[25]
port 100 nsew signal input
flabel metal3 s -800 5090 480 5202 0 FreeSans 1120 0 0 0 io_in_3v3[26]
port 101 nsew signal input
flabel metal3 s 583520 11000 584800 11112 0 FreeSans 1120 0 0 0 io_in_3v3[2]
port 102 nsew signal input
flabel metal3 s 583520 15728 584800 15840 0 FreeSans 1120 0 0 0 io_in_3v3[3]
port 103 nsew signal input
flabel metal3 s 583520 20456 584800 20568 0 FreeSans 1120 0 0 0 io_in_3v3[4]
port 104 nsew signal input
flabel metal3 s 583520 46914 584800 47026 0 FreeSans 1120 0 0 0 io_in_3v3[5]
port 105 nsew signal input
flabel metal3 s 583520 91572 584800 91684 0 FreeSans 1120 0 0 0 io_in_3v3[6]
port 106 nsew signal input
flabel metal3 s 583520 271594 584800 271706 0 FreeSans 1120 0 0 0 io_in_3v3[7]
port 107 nsew signal input
flabel metal3 s 583520 316016 584800 316128 0 FreeSans 1120 0 0 0 io_in_3v3[8]
port 108 nsew signal input
flabel metal3 s 583520 361238 584800 361350 0 FreeSans 1120 0 0 0 io_in_3v3[9]
port 109 nsew signal input
flabel metal3 s 583520 5090 584800 5202 0 FreeSans 1120 0 0 0 io_oeb[0]
port 110 nsew signal tristate
flabel metal3 s 583520 411206 584800 411318 0 FreeSans 1120 0 0 0 io_oeb[10]
port 111 nsew signal tristate
flabel metal3 s 583520 455628 584800 455740 0 FreeSans 1120 0 0 0 io_oeb[11]
port 112 nsew signal tristate
flabel metal3 s 583520 500050 584800 500162 0 FreeSans 1120 0 0 0 io_oeb[12]
port 113 nsew signal tristate
flabel metal3 s 583520 589472 584800 589584 0 FreeSans 1120 0 0 0 io_oeb[13]
port 114 nsew signal tristate
flabel metal3 s -800 505620 480 505732 0 FreeSans 1120 0 0 0 io_oeb[14]
port 115 nsew signal tristate
flabel metal3 s -800 462398 480 462510 0 FreeSans 1120 0 0 0 io_oeb[15]
port 116 nsew signal tristate
flabel metal3 s -800 419176 480 419288 0 FreeSans 1120 0 0 0 io_oeb[16]
port 117 nsew signal tristate
flabel metal3 s -800 375954 480 376066 0 FreeSans 1120 0 0 0 io_oeb[17]
port 118 nsew signal tristate
flabel metal3 s -800 332732 480 332844 0 FreeSans 1120 0 0 0 io_oeb[18]
port 119 nsew signal tristate
flabel metal3 s -800 289510 480 289622 0 FreeSans 1120 0 0 0 io_oeb[19]
port 120 nsew signal tristate
flabel metal3 s 583520 9818 584800 9930 0 FreeSans 1120 0 0 0 io_oeb[1]
port 121 nsew signal tristate
flabel metal3 s -800 246488 480 246600 0 FreeSans 1120 0 0 0 io_oeb[20]
port 122 nsew signal tristate
flabel metal3 s -800 118866 480 118978 0 FreeSans 1120 0 0 0 io_oeb[21]
port 123 nsew signal tristate
flabel metal3 s -800 75644 480 75756 0 FreeSans 1120 0 0 0 io_oeb[22]
port 124 nsew signal tristate
flabel metal3 s -800 32422 480 32534 0 FreeSans 1120 0 0 0 io_oeb[23]
port 125 nsew signal tristate
flabel metal3 s -800 11000 480 11112 0 FreeSans 1120 0 0 0 io_oeb[24]
port 126 nsew signal tristate
flabel metal3 s -800 6272 480 6384 0 FreeSans 1120 0 0 0 io_oeb[25]
port 127 nsew signal tristate
flabel metal3 s -800 1544 480 1656 0 FreeSans 1120 0 0 0 io_oeb[26]
port 128 nsew signal tristate
flabel metal3 s 583520 14546 584800 14658 0 FreeSans 1120 0 0 0 io_oeb[2]
port 129 nsew signal tristate
flabel metal3 s 583520 19274 584800 19386 0 FreeSans 1120 0 0 0 io_oeb[3]
port 130 nsew signal tristate
flabel metal3 s 583520 24002 584800 24114 0 FreeSans 1120 0 0 0 io_oeb[4]
port 131 nsew signal tristate
flabel metal3 s 583520 50460 584800 50572 0 FreeSans 1120 0 0 0 io_oeb[5]
port 132 nsew signal tristate
flabel metal3 s 583520 95118 584800 95230 0 FreeSans 1120 0 0 0 io_oeb[6]
port 133 nsew signal tristate
flabel metal3 s 583520 275140 584800 275252 0 FreeSans 1120 0 0 0 io_oeb[7]
port 134 nsew signal tristate
flabel metal3 s 583520 319562 584800 319674 0 FreeSans 1120 0 0 0 io_oeb[8]
port 135 nsew signal tristate
flabel metal3 s 583520 364784 584800 364896 0 FreeSans 1120 0 0 0 io_oeb[9]
port 136 nsew signal tristate
flabel metal3 s 583520 3908 584800 4020 0 FreeSans 1120 0 0 0 io_out[0]
port 137 nsew signal tristate
flabel metal3 s 583520 410024 584800 410136 0 FreeSans 1120 0 0 0 io_out[10]
port 138 nsew signal tristate
flabel metal3 s 583520 454446 584800 454558 0 FreeSans 1120 0 0 0 io_out[11]
port 139 nsew signal tristate
flabel metal3 s 583520 498868 584800 498980 0 FreeSans 1120 0 0 0 io_out[12]
port 140 nsew signal tristate
flabel metal3 s 583520 588290 584800 588402 0 FreeSans 1120 0 0 0 io_out[13]
port 141 nsew signal tristate
flabel metal3 s -800 506802 480 506914 0 FreeSans 1120 0 0 0 io_out[14]
port 142 nsew signal tristate
flabel metal3 s -800 463580 480 463692 0 FreeSans 1120 0 0 0 io_out[15]
port 143 nsew signal tristate
flabel metal3 s -800 420358 480 420470 0 FreeSans 1120 0 0 0 io_out[16]
port 144 nsew signal tristate
flabel metal3 s -800 377136 480 377248 0 FreeSans 1120 0 0 0 io_out[17]
port 145 nsew signal tristate
flabel metal3 s -800 333914 480 334026 0 FreeSans 1120 0 0 0 io_out[18]
port 146 nsew signal tristate
flabel metal3 s -800 290692 480 290804 0 FreeSans 1120 0 0 0 io_out[19]
port 147 nsew signal tristate
flabel metal3 s 583520 8636 584800 8748 0 FreeSans 1120 0 0 0 io_out[1]
port 148 nsew signal tristate
flabel metal3 s -800 247670 480 247782 0 FreeSans 1120 0 0 0 io_out[20]
port 149 nsew signal tristate
flabel metal3 s -800 120048 480 120160 0 FreeSans 1120 0 0 0 io_out[21]
port 150 nsew signal tristate
flabel metal3 s -800 76826 480 76938 0 FreeSans 1120 0 0 0 io_out[22]
port 151 nsew signal tristate
flabel metal3 s -800 33604 480 33716 0 FreeSans 1120 0 0 0 io_out[23]
port 152 nsew signal tristate
flabel metal3 s -800 12182 480 12294 0 FreeSans 1120 0 0 0 io_out[24]
port 153 nsew signal tristate
flabel metal3 s -800 7454 480 7566 0 FreeSans 1120 0 0 0 io_out[25]
port 154 nsew signal tristate
flabel metal3 s -800 2726 480 2838 0 FreeSans 1120 0 0 0 io_out[26]
port 155 nsew signal tristate
flabel metal3 s 583520 13364 584800 13476 0 FreeSans 1120 0 0 0 io_out[2]
port 156 nsew signal tristate
flabel metal3 s 583520 18092 584800 18204 0 FreeSans 1120 0 0 0 io_out[3]
port 157 nsew signal tristate
flabel metal3 s 583520 22820 584800 22932 0 FreeSans 1120 0 0 0 io_out[4]
port 158 nsew signal tristate
flabel metal3 s 583520 49278 584800 49390 0 FreeSans 1120 0 0 0 io_out[5]
port 159 nsew signal tristate
flabel metal3 s 583520 93936 584800 94048 0 FreeSans 1120 0 0 0 io_out[6]
port 160 nsew signal tristate
flabel metal3 s 583520 273958 584800 274070 0 FreeSans 1120 0 0 0 io_out[7]
port 161 nsew signal tristate
flabel metal3 s 583520 318380 584800 318492 0 FreeSans 1120 0 0 0 io_out[8]
port 162 nsew signal tristate
flabel metal3 s 583520 363602 584800 363714 0 FreeSans 1120 0 0 0 io_out[9]
port 163 nsew signal tristate
flabel metal2 s 125816 -800 125928 480 0 FreeSans 1120 90 0 0 la_data_in[0]
port 164 nsew signal input
flabel metal2 s 480416 -800 480528 480 0 FreeSans 1120 90 0 0 la_data_in[100]
port 165 nsew signal input
flabel metal2 s 483962 -800 484074 480 0 FreeSans 1120 90 0 0 la_data_in[101]
port 166 nsew signal input
flabel metal2 s 487508 -800 487620 480 0 FreeSans 1120 90 0 0 la_data_in[102]
port 167 nsew signal input
flabel metal2 s 491054 -800 491166 480 0 FreeSans 1120 90 0 0 la_data_in[103]
port 168 nsew signal input
flabel metal2 s 494600 -800 494712 480 0 FreeSans 1120 90 0 0 la_data_in[104]
port 169 nsew signal input
flabel metal2 s 498146 -800 498258 480 0 FreeSans 1120 90 0 0 la_data_in[105]
port 170 nsew signal input
flabel metal2 s 501692 -800 501804 480 0 FreeSans 1120 90 0 0 la_data_in[106]
port 171 nsew signal input
flabel metal2 s 505238 -800 505350 480 0 FreeSans 1120 90 0 0 la_data_in[107]
port 172 nsew signal input
flabel metal2 s 508784 -800 508896 480 0 FreeSans 1120 90 0 0 la_data_in[108]
port 173 nsew signal input
flabel metal2 s 512330 -800 512442 480 0 FreeSans 1120 90 0 0 la_data_in[109]
port 174 nsew signal input
flabel metal2 s 161276 -800 161388 480 0 FreeSans 1120 90 0 0 la_data_in[10]
port 175 nsew signal input
flabel metal2 s 515876 -800 515988 480 0 FreeSans 1120 90 0 0 la_data_in[110]
port 176 nsew signal input
flabel metal2 s 519422 -800 519534 480 0 FreeSans 1120 90 0 0 la_data_in[111]
port 177 nsew signal input
flabel metal2 s 522968 -800 523080 480 0 FreeSans 1120 90 0 0 la_data_in[112]
port 178 nsew signal input
flabel metal2 s 526514 -800 526626 480 0 FreeSans 1120 90 0 0 la_data_in[113]
port 179 nsew signal input
flabel metal2 s 530060 -800 530172 480 0 FreeSans 1120 90 0 0 la_data_in[114]
port 180 nsew signal input
flabel metal2 s 533606 -800 533718 480 0 FreeSans 1120 90 0 0 la_data_in[115]
port 181 nsew signal input
flabel metal2 s 537152 -800 537264 480 0 FreeSans 1120 90 0 0 la_data_in[116]
port 182 nsew signal input
flabel metal2 s 540698 -800 540810 480 0 FreeSans 1120 90 0 0 la_data_in[117]
port 183 nsew signal input
flabel metal2 s 544244 -800 544356 480 0 FreeSans 1120 90 0 0 la_data_in[118]
port 184 nsew signal input
flabel metal2 s 547790 -800 547902 480 0 FreeSans 1120 90 0 0 la_data_in[119]
port 185 nsew signal input
flabel metal2 s 164822 -800 164934 480 0 FreeSans 1120 90 0 0 la_data_in[11]
port 186 nsew signal input
flabel metal2 s 551336 -800 551448 480 0 FreeSans 1120 90 0 0 la_data_in[120]
port 187 nsew signal input
flabel metal2 s 554882 -800 554994 480 0 FreeSans 1120 90 0 0 la_data_in[121]
port 188 nsew signal input
flabel metal2 s 558428 -800 558540 480 0 FreeSans 1120 90 0 0 la_data_in[122]
port 189 nsew signal input
flabel metal2 s 561974 -800 562086 480 0 FreeSans 1120 90 0 0 la_data_in[123]
port 190 nsew signal input
flabel metal2 s 565520 -800 565632 480 0 FreeSans 1120 90 0 0 la_data_in[124]
port 191 nsew signal input
flabel metal2 s 569066 -800 569178 480 0 FreeSans 1120 90 0 0 la_data_in[125]
port 192 nsew signal input
flabel metal2 s 572612 -800 572724 480 0 FreeSans 1120 90 0 0 la_data_in[126]
port 193 nsew signal input
flabel metal2 s 576158 -800 576270 480 0 FreeSans 1120 90 0 0 la_data_in[127]
port 194 nsew signal input
flabel metal2 s 168368 -800 168480 480 0 FreeSans 1120 90 0 0 la_data_in[12]
port 195 nsew signal input
flabel metal2 s 171914 -800 172026 480 0 FreeSans 1120 90 0 0 la_data_in[13]
port 196 nsew signal input
flabel metal2 s 175460 -800 175572 480 0 FreeSans 1120 90 0 0 la_data_in[14]
port 197 nsew signal input
flabel metal2 s 179006 -800 179118 480 0 FreeSans 1120 90 0 0 la_data_in[15]
port 198 nsew signal input
flabel metal2 s 182552 -800 182664 480 0 FreeSans 1120 90 0 0 la_data_in[16]
port 199 nsew signal input
flabel metal2 s 186098 -800 186210 480 0 FreeSans 1120 90 0 0 la_data_in[17]
port 200 nsew signal input
flabel metal2 s 189644 -800 189756 480 0 FreeSans 1120 90 0 0 la_data_in[18]
port 201 nsew signal input
flabel metal2 s 193190 -800 193302 480 0 FreeSans 1120 90 0 0 la_data_in[19]
port 202 nsew signal input
flabel metal2 s 129362 -800 129474 480 0 FreeSans 1120 90 0 0 la_data_in[1]
port 203 nsew signal input
flabel metal2 s 196736 -800 196848 480 0 FreeSans 1120 90 0 0 la_data_in[20]
port 204 nsew signal input
flabel metal2 s 200282 -800 200394 480 0 FreeSans 1120 90 0 0 la_data_in[21]
port 205 nsew signal input
flabel metal2 s 203828 -800 203940 480 0 FreeSans 1120 90 0 0 la_data_in[22]
port 206 nsew signal input
flabel metal2 s 207374 -800 207486 480 0 FreeSans 1120 90 0 0 la_data_in[23]
port 207 nsew signal input
flabel metal2 s 210920 -800 211032 480 0 FreeSans 1120 90 0 0 la_data_in[24]
port 208 nsew signal input
flabel metal2 s 214466 -800 214578 480 0 FreeSans 1120 90 0 0 la_data_in[25]
port 209 nsew signal input
flabel metal2 s 218012 -800 218124 480 0 FreeSans 1120 90 0 0 la_data_in[26]
port 210 nsew signal input
flabel metal2 s 221558 -800 221670 480 0 FreeSans 1120 90 0 0 la_data_in[27]
port 211 nsew signal input
flabel metal2 s 225104 -800 225216 480 0 FreeSans 1120 90 0 0 la_data_in[28]
port 212 nsew signal input
flabel metal2 s 228650 -800 228762 480 0 FreeSans 1120 90 0 0 la_data_in[29]
port 213 nsew signal input
flabel metal2 s 132908 -800 133020 480 0 FreeSans 1120 90 0 0 la_data_in[2]
port 214 nsew signal input
flabel metal2 s 232196 -800 232308 480 0 FreeSans 1120 90 0 0 la_data_in[30]
port 215 nsew signal input
flabel metal2 s 235742 -800 235854 480 0 FreeSans 1120 90 0 0 la_data_in[31]
port 216 nsew signal input
flabel metal2 s 239288 -800 239400 480 0 FreeSans 1120 90 0 0 la_data_in[32]
port 217 nsew signal input
flabel metal2 s 242834 -800 242946 480 0 FreeSans 1120 90 0 0 la_data_in[33]
port 218 nsew signal input
flabel metal2 s 246380 -800 246492 480 0 FreeSans 1120 90 0 0 la_data_in[34]
port 219 nsew signal input
flabel metal2 s 249926 -800 250038 480 0 FreeSans 1120 90 0 0 la_data_in[35]
port 220 nsew signal input
flabel metal2 s 253472 -800 253584 480 0 FreeSans 1120 90 0 0 la_data_in[36]
port 221 nsew signal input
flabel metal2 s 257018 -800 257130 480 0 FreeSans 1120 90 0 0 la_data_in[37]
port 222 nsew signal input
flabel metal2 s 260564 -800 260676 480 0 FreeSans 1120 90 0 0 la_data_in[38]
port 223 nsew signal input
flabel metal2 s 264110 -800 264222 480 0 FreeSans 1120 90 0 0 la_data_in[39]
port 224 nsew signal input
flabel metal2 s 136454 -800 136566 480 0 FreeSans 1120 90 0 0 la_data_in[3]
port 225 nsew signal input
flabel metal2 s 267656 -800 267768 480 0 FreeSans 1120 90 0 0 la_data_in[40]
port 226 nsew signal input
flabel metal2 s 271202 -800 271314 480 0 FreeSans 1120 90 0 0 la_data_in[41]
port 227 nsew signal input
flabel metal2 s 274748 -800 274860 480 0 FreeSans 1120 90 0 0 la_data_in[42]
port 228 nsew signal input
flabel metal2 s 278294 -800 278406 480 0 FreeSans 1120 90 0 0 la_data_in[43]
port 229 nsew signal input
flabel metal2 s 281840 -800 281952 480 0 FreeSans 1120 90 0 0 la_data_in[44]
port 230 nsew signal input
flabel metal2 s 285386 -800 285498 480 0 FreeSans 1120 90 0 0 la_data_in[45]
port 231 nsew signal input
flabel metal2 s 288932 -800 289044 480 0 FreeSans 1120 90 0 0 la_data_in[46]
port 232 nsew signal input
flabel metal2 s 292478 -800 292590 480 0 FreeSans 1120 90 0 0 la_data_in[47]
port 233 nsew signal input
flabel metal2 s 296024 -800 296136 480 0 FreeSans 1120 90 0 0 la_data_in[48]
port 234 nsew signal input
flabel metal2 s 299570 -800 299682 480 0 FreeSans 1120 90 0 0 la_data_in[49]
port 235 nsew signal input
flabel metal2 s 140000 -800 140112 480 0 FreeSans 1120 90 0 0 la_data_in[4]
port 236 nsew signal input
flabel metal2 s 303116 -800 303228 480 0 FreeSans 1120 90 0 0 la_data_in[50]
port 237 nsew signal input
flabel metal2 s 306662 -800 306774 480 0 FreeSans 1120 90 0 0 la_data_in[51]
port 238 nsew signal input
flabel metal2 s 310208 -800 310320 480 0 FreeSans 1120 90 0 0 la_data_in[52]
port 239 nsew signal input
flabel metal2 s 313754 -800 313866 480 0 FreeSans 1120 90 0 0 la_data_in[53]
port 240 nsew signal input
flabel metal2 s 317300 -800 317412 480 0 FreeSans 1120 90 0 0 la_data_in[54]
port 241 nsew signal input
flabel metal2 s 320846 -800 320958 480 0 FreeSans 1120 90 0 0 la_data_in[55]
port 242 nsew signal input
flabel metal2 s 324392 -800 324504 480 0 FreeSans 1120 90 0 0 la_data_in[56]
port 243 nsew signal input
flabel metal2 s 327938 -800 328050 480 0 FreeSans 1120 90 0 0 la_data_in[57]
port 244 nsew signal input
flabel metal2 s 331484 -800 331596 480 0 FreeSans 1120 90 0 0 la_data_in[58]
port 245 nsew signal input
flabel metal2 s 335030 -800 335142 480 0 FreeSans 1120 90 0 0 la_data_in[59]
port 246 nsew signal input
flabel metal2 s 143546 -800 143658 480 0 FreeSans 1120 90 0 0 la_data_in[5]
port 247 nsew signal input
flabel metal2 s 338576 -800 338688 480 0 FreeSans 1120 90 0 0 la_data_in[60]
port 248 nsew signal input
flabel metal2 s 342122 -800 342234 480 0 FreeSans 1120 90 0 0 la_data_in[61]
port 249 nsew signal input
flabel metal2 s 345668 -800 345780 480 0 FreeSans 1120 90 0 0 la_data_in[62]
port 250 nsew signal input
flabel metal2 s 349214 -800 349326 480 0 FreeSans 1120 90 0 0 la_data_in[63]
port 251 nsew signal input
flabel metal2 s 352760 -800 352872 480 0 FreeSans 1120 90 0 0 la_data_in[64]
port 252 nsew signal input
flabel metal2 s 356306 -800 356418 480 0 FreeSans 1120 90 0 0 la_data_in[65]
port 253 nsew signal input
flabel metal2 s 359852 -800 359964 480 0 FreeSans 1120 90 0 0 la_data_in[66]
port 254 nsew signal input
flabel metal2 s 363398 -800 363510 480 0 FreeSans 1120 90 0 0 la_data_in[67]
port 255 nsew signal input
flabel metal2 s 366944 -800 367056 480 0 FreeSans 1120 90 0 0 la_data_in[68]
port 256 nsew signal input
flabel metal2 s 370490 -800 370602 480 0 FreeSans 1120 90 0 0 la_data_in[69]
port 257 nsew signal input
flabel metal2 s 147092 -800 147204 480 0 FreeSans 1120 90 0 0 la_data_in[6]
port 258 nsew signal input
flabel metal2 s 374036 -800 374148 480 0 FreeSans 1120 90 0 0 la_data_in[70]
port 259 nsew signal input
flabel metal2 s 377582 -800 377694 480 0 FreeSans 1120 90 0 0 la_data_in[71]
port 260 nsew signal input
flabel metal2 s 381128 -800 381240 480 0 FreeSans 1120 90 0 0 la_data_in[72]
port 261 nsew signal input
flabel metal2 s 384674 -800 384786 480 0 FreeSans 1120 90 0 0 la_data_in[73]
port 262 nsew signal input
flabel metal2 s 388220 -800 388332 480 0 FreeSans 1120 90 0 0 la_data_in[74]
port 263 nsew signal input
flabel metal2 s 391766 -800 391878 480 0 FreeSans 1120 90 0 0 la_data_in[75]
port 264 nsew signal input
flabel metal2 s 395312 -800 395424 480 0 FreeSans 1120 90 0 0 la_data_in[76]
port 265 nsew signal input
flabel metal2 s 398858 -800 398970 480 0 FreeSans 1120 90 0 0 la_data_in[77]
port 266 nsew signal input
flabel metal2 s 402404 -800 402516 480 0 FreeSans 1120 90 0 0 la_data_in[78]
port 267 nsew signal input
flabel metal2 s 405950 -800 406062 480 0 FreeSans 1120 90 0 0 la_data_in[79]
port 268 nsew signal input
flabel metal2 s 150638 -800 150750 480 0 FreeSans 1120 90 0 0 la_data_in[7]
port 269 nsew signal input
flabel metal2 s 409496 -800 409608 480 0 FreeSans 1120 90 0 0 la_data_in[80]
port 270 nsew signal input
flabel metal2 s 413042 -800 413154 480 0 FreeSans 1120 90 0 0 la_data_in[81]
port 271 nsew signal input
flabel metal2 s 416588 -800 416700 480 0 FreeSans 1120 90 0 0 la_data_in[82]
port 272 nsew signal input
flabel metal2 s 420134 -800 420246 480 0 FreeSans 1120 90 0 0 la_data_in[83]
port 273 nsew signal input
flabel metal2 s 423680 -800 423792 480 0 FreeSans 1120 90 0 0 la_data_in[84]
port 274 nsew signal input
flabel metal2 s 427226 -800 427338 480 0 FreeSans 1120 90 0 0 la_data_in[85]
port 275 nsew signal input
flabel metal2 s 430772 -800 430884 480 0 FreeSans 1120 90 0 0 la_data_in[86]
port 276 nsew signal input
flabel metal2 s 434318 -800 434430 480 0 FreeSans 1120 90 0 0 la_data_in[87]
port 277 nsew signal input
flabel metal2 s 437864 -800 437976 480 0 FreeSans 1120 90 0 0 la_data_in[88]
port 278 nsew signal input
flabel metal2 s 441410 -800 441522 480 0 FreeSans 1120 90 0 0 la_data_in[89]
port 279 nsew signal input
flabel metal2 s 154184 -800 154296 480 0 FreeSans 1120 90 0 0 la_data_in[8]
port 280 nsew signal input
flabel metal2 s 444956 -800 445068 480 0 FreeSans 1120 90 0 0 la_data_in[90]
port 281 nsew signal input
flabel metal2 s 448502 -800 448614 480 0 FreeSans 1120 90 0 0 la_data_in[91]
port 282 nsew signal input
flabel metal2 s 452048 -800 452160 480 0 FreeSans 1120 90 0 0 la_data_in[92]
port 283 nsew signal input
flabel metal2 s 455594 -800 455706 480 0 FreeSans 1120 90 0 0 la_data_in[93]
port 284 nsew signal input
flabel metal2 s 459140 -800 459252 480 0 FreeSans 1120 90 0 0 la_data_in[94]
port 285 nsew signal input
flabel metal2 s 462686 -800 462798 480 0 FreeSans 1120 90 0 0 la_data_in[95]
port 286 nsew signal input
flabel metal2 s 466232 -800 466344 480 0 FreeSans 1120 90 0 0 la_data_in[96]
port 287 nsew signal input
flabel metal2 s 469778 -800 469890 480 0 FreeSans 1120 90 0 0 la_data_in[97]
port 288 nsew signal input
flabel metal2 s 473324 -800 473436 480 0 FreeSans 1120 90 0 0 la_data_in[98]
port 289 nsew signal input
flabel metal2 s 476870 -800 476982 480 0 FreeSans 1120 90 0 0 la_data_in[99]
port 290 nsew signal input
flabel metal2 s 157730 -800 157842 480 0 FreeSans 1120 90 0 0 la_data_in[9]
port 291 nsew signal input
flabel metal2 s 126998 -800 127110 480 0 FreeSans 1120 90 0 0 la_data_out[0]
port 292 nsew signal tristate
flabel metal2 s 481598 -800 481710 480 0 FreeSans 1120 90 0 0 la_data_out[100]
port 293 nsew signal tristate
flabel metal2 s 485144 -800 485256 480 0 FreeSans 1120 90 0 0 la_data_out[101]
port 294 nsew signal tristate
flabel metal2 s 488690 -800 488802 480 0 FreeSans 1120 90 0 0 la_data_out[102]
port 295 nsew signal tristate
flabel metal2 s 492236 -800 492348 480 0 FreeSans 1120 90 0 0 la_data_out[103]
port 296 nsew signal tristate
flabel metal2 s 495782 -800 495894 480 0 FreeSans 1120 90 0 0 la_data_out[104]
port 297 nsew signal tristate
flabel metal2 s 499328 -800 499440 480 0 FreeSans 1120 90 0 0 la_data_out[105]
port 298 nsew signal tristate
flabel metal2 s 502874 -800 502986 480 0 FreeSans 1120 90 0 0 la_data_out[106]
port 299 nsew signal tristate
flabel metal2 s 506420 -800 506532 480 0 FreeSans 1120 90 0 0 la_data_out[107]
port 300 nsew signal tristate
flabel metal2 s 509966 -800 510078 480 0 FreeSans 1120 90 0 0 la_data_out[108]
port 301 nsew signal tristate
flabel metal2 s 513512 -800 513624 480 0 FreeSans 1120 90 0 0 la_data_out[109]
port 302 nsew signal tristate
flabel metal2 s 162458 -800 162570 480 0 FreeSans 1120 90 0 0 la_data_out[10]
port 303 nsew signal tristate
flabel metal2 s 517058 -800 517170 480 0 FreeSans 1120 90 0 0 la_data_out[110]
port 304 nsew signal tristate
flabel metal2 s 520604 -800 520716 480 0 FreeSans 1120 90 0 0 la_data_out[111]
port 305 nsew signal tristate
flabel metal2 s 524150 -800 524262 480 0 FreeSans 1120 90 0 0 la_data_out[112]
port 306 nsew signal tristate
flabel metal2 s 527696 -800 527808 480 0 FreeSans 1120 90 0 0 la_data_out[113]
port 307 nsew signal tristate
flabel metal2 s 531242 -800 531354 480 0 FreeSans 1120 90 0 0 la_data_out[114]
port 308 nsew signal tristate
flabel metal2 s 534788 -800 534900 480 0 FreeSans 1120 90 0 0 la_data_out[115]
port 309 nsew signal tristate
flabel metal2 s 538334 -800 538446 480 0 FreeSans 1120 90 0 0 la_data_out[116]
port 310 nsew signal tristate
flabel metal2 s 541880 -800 541992 480 0 FreeSans 1120 90 0 0 la_data_out[117]
port 311 nsew signal tristate
flabel metal2 s 545426 -800 545538 480 0 FreeSans 1120 90 0 0 la_data_out[118]
port 312 nsew signal tristate
flabel metal2 s 548972 -800 549084 480 0 FreeSans 1120 90 0 0 la_data_out[119]
port 313 nsew signal tristate
flabel metal2 s 166004 -800 166116 480 0 FreeSans 1120 90 0 0 la_data_out[11]
port 314 nsew signal tristate
flabel metal2 s 552518 -800 552630 480 0 FreeSans 1120 90 0 0 la_data_out[120]
port 315 nsew signal tristate
flabel metal2 s 556064 -800 556176 480 0 FreeSans 1120 90 0 0 la_data_out[121]
port 316 nsew signal tristate
flabel metal2 s 559610 -800 559722 480 0 FreeSans 1120 90 0 0 la_data_out[122]
port 317 nsew signal tristate
flabel metal2 s 563156 -800 563268 480 0 FreeSans 1120 90 0 0 la_data_out[123]
port 318 nsew signal tristate
flabel metal2 s 566702 -800 566814 480 0 FreeSans 1120 90 0 0 la_data_out[124]
port 319 nsew signal tristate
flabel metal2 s 570248 -800 570360 480 0 FreeSans 1120 90 0 0 la_data_out[125]
port 320 nsew signal tristate
flabel metal2 s 573794 -800 573906 480 0 FreeSans 1120 90 0 0 la_data_out[126]
port 321 nsew signal tristate
flabel metal2 s 577340 -800 577452 480 0 FreeSans 1120 90 0 0 la_data_out[127]
port 322 nsew signal tristate
flabel metal2 s 169550 -800 169662 480 0 FreeSans 1120 90 0 0 la_data_out[12]
port 323 nsew signal tristate
flabel metal2 s 173096 -800 173208 480 0 FreeSans 1120 90 0 0 la_data_out[13]
port 324 nsew signal tristate
flabel metal2 s 176642 -800 176754 480 0 FreeSans 1120 90 0 0 la_data_out[14]
port 325 nsew signal tristate
flabel metal2 s 180188 -800 180300 480 0 FreeSans 1120 90 0 0 la_data_out[15]
port 326 nsew signal tristate
flabel metal2 s 183734 -800 183846 480 0 FreeSans 1120 90 0 0 la_data_out[16]
port 327 nsew signal tristate
flabel metal2 s 187280 -800 187392 480 0 FreeSans 1120 90 0 0 la_data_out[17]
port 328 nsew signal tristate
flabel metal2 s 190826 -800 190938 480 0 FreeSans 1120 90 0 0 la_data_out[18]
port 329 nsew signal tristate
flabel metal2 s 194372 -800 194484 480 0 FreeSans 1120 90 0 0 la_data_out[19]
port 330 nsew signal tristate
flabel metal2 s 130544 -800 130656 480 0 FreeSans 1120 90 0 0 la_data_out[1]
port 331 nsew signal tristate
flabel metal2 s 197918 -800 198030 480 0 FreeSans 1120 90 0 0 la_data_out[20]
port 332 nsew signal tristate
flabel metal2 s 201464 -800 201576 480 0 FreeSans 1120 90 0 0 la_data_out[21]
port 333 nsew signal tristate
flabel metal2 s 205010 -800 205122 480 0 FreeSans 1120 90 0 0 la_data_out[22]
port 334 nsew signal tristate
flabel metal2 s 208556 -800 208668 480 0 FreeSans 1120 90 0 0 la_data_out[23]
port 335 nsew signal tristate
flabel metal2 s 212102 -800 212214 480 0 FreeSans 1120 90 0 0 la_data_out[24]
port 336 nsew signal tristate
flabel metal2 s 215648 -800 215760 480 0 FreeSans 1120 90 0 0 la_data_out[25]
port 337 nsew signal tristate
flabel metal2 s 219194 -800 219306 480 0 FreeSans 1120 90 0 0 la_data_out[26]
port 338 nsew signal tristate
flabel metal2 s 222740 -800 222852 480 0 FreeSans 1120 90 0 0 la_data_out[27]
port 339 nsew signal tristate
flabel metal2 s 226286 -800 226398 480 0 FreeSans 1120 90 0 0 la_data_out[28]
port 340 nsew signal tristate
flabel metal2 s 229832 -800 229944 480 0 FreeSans 1120 90 0 0 la_data_out[29]
port 341 nsew signal tristate
flabel metal2 s 134090 -800 134202 480 0 FreeSans 1120 90 0 0 la_data_out[2]
port 342 nsew signal tristate
flabel metal2 s 233378 -800 233490 480 0 FreeSans 1120 90 0 0 la_data_out[30]
port 343 nsew signal tristate
flabel metal2 s 236924 -800 237036 480 0 FreeSans 1120 90 0 0 la_data_out[31]
port 344 nsew signal tristate
flabel metal2 s 240470 -800 240582 480 0 FreeSans 1120 90 0 0 la_data_out[32]
port 345 nsew signal tristate
flabel metal2 s 244016 -800 244128 480 0 FreeSans 1120 90 0 0 la_data_out[33]
port 346 nsew signal tristate
flabel metal2 s 247562 -800 247674 480 0 FreeSans 1120 90 0 0 la_data_out[34]
port 347 nsew signal tristate
flabel metal2 s 251108 -800 251220 480 0 FreeSans 1120 90 0 0 la_data_out[35]
port 348 nsew signal tristate
flabel metal2 s 254654 -800 254766 480 0 FreeSans 1120 90 0 0 la_data_out[36]
port 349 nsew signal tristate
flabel metal2 s 258200 -800 258312 480 0 FreeSans 1120 90 0 0 la_data_out[37]
port 350 nsew signal tristate
flabel metal2 s 261746 -800 261858 480 0 FreeSans 1120 90 0 0 la_data_out[38]
port 351 nsew signal tristate
flabel metal2 s 265292 -800 265404 480 0 FreeSans 1120 90 0 0 la_data_out[39]
port 352 nsew signal tristate
flabel metal2 s 137636 -800 137748 480 0 FreeSans 1120 90 0 0 la_data_out[3]
port 353 nsew signal tristate
flabel metal2 s 268838 -800 268950 480 0 FreeSans 1120 90 0 0 la_data_out[40]
port 354 nsew signal tristate
flabel metal2 s 272384 -800 272496 480 0 FreeSans 1120 90 0 0 la_data_out[41]
port 355 nsew signal tristate
flabel metal2 s 275930 -800 276042 480 0 FreeSans 1120 90 0 0 la_data_out[42]
port 356 nsew signal tristate
flabel metal2 s 279476 -800 279588 480 0 FreeSans 1120 90 0 0 la_data_out[43]
port 357 nsew signal tristate
flabel metal2 s 283022 -800 283134 480 0 FreeSans 1120 90 0 0 la_data_out[44]
port 358 nsew signal tristate
flabel metal2 s 286568 -800 286680 480 0 FreeSans 1120 90 0 0 la_data_out[45]
port 359 nsew signal tristate
flabel metal2 s 290114 -800 290226 480 0 FreeSans 1120 90 0 0 la_data_out[46]
port 360 nsew signal tristate
flabel metal2 s 293660 -800 293772 480 0 FreeSans 1120 90 0 0 la_data_out[47]
port 361 nsew signal tristate
flabel metal2 s 297206 -800 297318 480 0 FreeSans 1120 90 0 0 la_data_out[48]
port 362 nsew signal tristate
flabel metal2 s 300752 -800 300864 480 0 FreeSans 1120 90 0 0 la_data_out[49]
port 363 nsew signal tristate
flabel metal2 s 141182 -800 141294 480 0 FreeSans 1120 90 0 0 la_data_out[4]
port 364 nsew signal tristate
flabel metal2 s 304298 -800 304410 480 0 FreeSans 1120 90 0 0 la_data_out[50]
port 365 nsew signal tristate
flabel metal2 s 307844 -800 307956 480 0 FreeSans 1120 90 0 0 la_data_out[51]
port 366 nsew signal tristate
flabel metal2 s 311390 -800 311502 480 0 FreeSans 1120 90 0 0 la_data_out[52]
port 367 nsew signal tristate
flabel metal2 s 314936 -800 315048 480 0 FreeSans 1120 90 0 0 la_data_out[53]
port 368 nsew signal tristate
flabel metal2 s 318482 -800 318594 480 0 FreeSans 1120 90 0 0 la_data_out[54]
port 369 nsew signal tristate
flabel metal2 s 322028 -800 322140 480 0 FreeSans 1120 90 0 0 la_data_out[55]
port 370 nsew signal tristate
flabel metal2 s 325574 -800 325686 480 0 FreeSans 1120 90 0 0 la_data_out[56]
port 371 nsew signal tristate
flabel metal2 s 329120 -800 329232 480 0 FreeSans 1120 90 0 0 la_data_out[57]
port 372 nsew signal tristate
flabel metal2 s 332666 -800 332778 480 0 FreeSans 1120 90 0 0 la_data_out[58]
port 373 nsew signal tristate
flabel metal2 s 336212 -800 336324 480 0 FreeSans 1120 90 0 0 la_data_out[59]
port 374 nsew signal tristate
flabel metal2 s 144728 -800 144840 480 0 FreeSans 1120 90 0 0 la_data_out[5]
port 375 nsew signal tristate
flabel metal2 s 339758 -800 339870 480 0 FreeSans 1120 90 0 0 la_data_out[60]
port 376 nsew signal tristate
flabel metal2 s 343304 -800 343416 480 0 FreeSans 1120 90 0 0 la_data_out[61]
port 377 nsew signal tristate
flabel metal2 s 346850 -800 346962 480 0 FreeSans 1120 90 0 0 la_data_out[62]
port 378 nsew signal tristate
flabel metal2 s 350396 -800 350508 480 0 FreeSans 1120 90 0 0 la_data_out[63]
port 379 nsew signal tristate
flabel metal2 s 353942 -800 354054 480 0 FreeSans 1120 90 0 0 la_data_out[64]
port 380 nsew signal tristate
flabel metal2 s 357488 -800 357600 480 0 FreeSans 1120 90 0 0 la_data_out[65]
port 381 nsew signal tristate
flabel metal2 s 361034 -800 361146 480 0 FreeSans 1120 90 0 0 la_data_out[66]
port 382 nsew signal tristate
flabel metal2 s 364580 -800 364692 480 0 FreeSans 1120 90 0 0 la_data_out[67]
port 383 nsew signal tristate
flabel metal2 s 368126 -800 368238 480 0 FreeSans 1120 90 0 0 la_data_out[68]
port 384 nsew signal tristate
flabel metal2 s 371672 -800 371784 480 0 FreeSans 1120 90 0 0 la_data_out[69]
port 385 nsew signal tristate
flabel metal2 s 148274 -800 148386 480 0 FreeSans 1120 90 0 0 la_data_out[6]
port 386 nsew signal tristate
flabel metal2 s 375218 -800 375330 480 0 FreeSans 1120 90 0 0 la_data_out[70]
port 387 nsew signal tristate
flabel metal2 s 378764 -800 378876 480 0 FreeSans 1120 90 0 0 la_data_out[71]
port 388 nsew signal tristate
flabel metal2 s 382310 -800 382422 480 0 FreeSans 1120 90 0 0 la_data_out[72]
port 389 nsew signal tristate
flabel metal2 s 385856 -800 385968 480 0 FreeSans 1120 90 0 0 la_data_out[73]
port 390 nsew signal tristate
flabel metal2 s 389402 -800 389514 480 0 FreeSans 1120 90 0 0 la_data_out[74]
port 391 nsew signal tristate
flabel metal2 s 392948 -800 393060 480 0 FreeSans 1120 90 0 0 la_data_out[75]
port 392 nsew signal tristate
flabel metal2 s 396494 -800 396606 480 0 FreeSans 1120 90 0 0 la_data_out[76]
port 393 nsew signal tristate
flabel metal2 s 400040 -800 400152 480 0 FreeSans 1120 90 0 0 la_data_out[77]
port 394 nsew signal tristate
flabel metal2 s 403586 -800 403698 480 0 FreeSans 1120 90 0 0 la_data_out[78]
port 395 nsew signal tristate
flabel metal2 s 407132 -800 407244 480 0 FreeSans 1120 90 0 0 la_data_out[79]
port 396 nsew signal tristate
flabel metal2 s 151820 -800 151932 480 0 FreeSans 1120 90 0 0 la_data_out[7]
port 397 nsew signal tristate
flabel metal2 s 410678 -800 410790 480 0 FreeSans 1120 90 0 0 la_data_out[80]
port 398 nsew signal tristate
flabel metal2 s 414224 -800 414336 480 0 FreeSans 1120 90 0 0 la_data_out[81]
port 399 nsew signal tristate
flabel metal2 s 417770 -800 417882 480 0 FreeSans 1120 90 0 0 la_data_out[82]
port 400 nsew signal tristate
flabel metal2 s 421316 -800 421428 480 0 FreeSans 1120 90 0 0 la_data_out[83]
port 401 nsew signal tristate
flabel metal2 s 424862 -800 424974 480 0 FreeSans 1120 90 0 0 la_data_out[84]
port 402 nsew signal tristate
flabel metal2 s 428408 -800 428520 480 0 FreeSans 1120 90 0 0 la_data_out[85]
port 403 nsew signal tristate
flabel metal2 s 431954 -800 432066 480 0 FreeSans 1120 90 0 0 la_data_out[86]
port 404 nsew signal tristate
flabel metal2 s 435500 -800 435612 480 0 FreeSans 1120 90 0 0 la_data_out[87]
port 405 nsew signal tristate
flabel metal2 s 439046 -800 439158 480 0 FreeSans 1120 90 0 0 la_data_out[88]
port 406 nsew signal tristate
flabel metal2 s 442592 -800 442704 480 0 FreeSans 1120 90 0 0 la_data_out[89]
port 407 nsew signal tristate
flabel metal2 s 155366 -800 155478 480 0 FreeSans 1120 90 0 0 la_data_out[8]
port 408 nsew signal tristate
flabel metal2 s 446138 -800 446250 480 0 FreeSans 1120 90 0 0 la_data_out[90]
port 409 nsew signal tristate
flabel metal2 s 449684 -800 449796 480 0 FreeSans 1120 90 0 0 la_data_out[91]
port 410 nsew signal tristate
flabel metal2 s 453230 -800 453342 480 0 FreeSans 1120 90 0 0 la_data_out[92]
port 411 nsew signal tristate
flabel metal2 s 456776 -800 456888 480 0 FreeSans 1120 90 0 0 la_data_out[93]
port 412 nsew signal tristate
flabel metal2 s 460322 -800 460434 480 0 FreeSans 1120 90 0 0 la_data_out[94]
port 413 nsew signal tristate
flabel metal2 s 463868 -800 463980 480 0 FreeSans 1120 90 0 0 la_data_out[95]
port 414 nsew signal tristate
flabel metal2 s 467414 -800 467526 480 0 FreeSans 1120 90 0 0 la_data_out[96]
port 415 nsew signal tristate
flabel metal2 s 470960 -800 471072 480 0 FreeSans 1120 90 0 0 la_data_out[97]
port 416 nsew signal tristate
flabel metal2 s 474506 -800 474618 480 0 FreeSans 1120 90 0 0 la_data_out[98]
port 417 nsew signal tristate
flabel metal2 s 478052 -800 478164 480 0 FreeSans 1120 90 0 0 la_data_out[99]
port 418 nsew signal tristate
flabel metal2 s 158912 -800 159024 480 0 FreeSans 1120 90 0 0 la_data_out[9]
port 419 nsew signal tristate
flabel metal2 s 128180 -800 128292 480 0 FreeSans 1120 90 0 0 la_oenb[0]
port 420 nsew signal input
flabel metal2 s 482780 -800 482892 480 0 FreeSans 1120 90 0 0 la_oenb[100]
port 421 nsew signal input
flabel metal2 s 486326 -800 486438 480 0 FreeSans 1120 90 0 0 la_oenb[101]
port 422 nsew signal input
flabel metal2 s 489872 -800 489984 480 0 FreeSans 1120 90 0 0 la_oenb[102]
port 423 nsew signal input
flabel metal2 s 493418 -800 493530 480 0 FreeSans 1120 90 0 0 la_oenb[103]
port 424 nsew signal input
flabel metal2 s 496964 -800 497076 480 0 FreeSans 1120 90 0 0 la_oenb[104]
port 425 nsew signal input
flabel metal2 s 500510 -800 500622 480 0 FreeSans 1120 90 0 0 la_oenb[105]
port 426 nsew signal input
flabel metal2 s 504056 -800 504168 480 0 FreeSans 1120 90 0 0 la_oenb[106]
port 427 nsew signal input
flabel metal2 s 507602 -800 507714 480 0 FreeSans 1120 90 0 0 la_oenb[107]
port 428 nsew signal input
flabel metal2 s 511148 -800 511260 480 0 FreeSans 1120 90 0 0 la_oenb[108]
port 429 nsew signal input
flabel metal2 s 514694 -800 514806 480 0 FreeSans 1120 90 0 0 la_oenb[109]
port 430 nsew signal input
flabel metal2 s 163640 -800 163752 480 0 FreeSans 1120 90 0 0 la_oenb[10]
port 431 nsew signal input
flabel metal2 s 518240 -800 518352 480 0 FreeSans 1120 90 0 0 la_oenb[110]
port 432 nsew signal input
flabel metal2 s 521786 -800 521898 480 0 FreeSans 1120 90 0 0 la_oenb[111]
port 433 nsew signal input
flabel metal2 s 525332 -800 525444 480 0 FreeSans 1120 90 0 0 la_oenb[112]
port 434 nsew signal input
flabel metal2 s 528878 -800 528990 480 0 FreeSans 1120 90 0 0 la_oenb[113]
port 435 nsew signal input
flabel metal2 s 532424 -800 532536 480 0 FreeSans 1120 90 0 0 la_oenb[114]
port 436 nsew signal input
flabel metal2 s 535970 -800 536082 480 0 FreeSans 1120 90 0 0 la_oenb[115]
port 437 nsew signal input
flabel metal2 s 539516 -800 539628 480 0 FreeSans 1120 90 0 0 la_oenb[116]
port 438 nsew signal input
flabel metal2 s 543062 -800 543174 480 0 FreeSans 1120 90 0 0 la_oenb[117]
port 439 nsew signal input
flabel metal2 s 546608 -800 546720 480 0 FreeSans 1120 90 0 0 la_oenb[118]
port 440 nsew signal input
flabel metal2 s 550154 -800 550266 480 0 FreeSans 1120 90 0 0 la_oenb[119]
port 441 nsew signal input
flabel metal2 s 167186 -800 167298 480 0 FreeSans 1120 90 0 0 la_oenb[11]
port 442 nsew signal input
flabel metal2 s 553700 -800 553812 480 0 FreeSans 1120 90 0 0 la_oenb[120]
port 443 nsew signal input
flabel metal2 s 557246 -800 557358 480 0 FreeSans 1120 90 0 0 la_oenb[121]
port 444 nsew signal input
flabel metal2 s 560792 -800 560904 480 0 FreeSans 1120 90 0 0 la_oenb[122]
port 445 nsew signal input
flabel metal2 s 564338 -800 564450 480 0 FreeSans 1120 90 0 0 la_oenb[123]
port 446 nsew signal input
flabel metal2 s 567884 -800 567996 480 0 FreeSans 1120 90 0 0 la_oenb[124]
port 447 nsew signal input
flabel metal2 s 571430 -800 571542 480 0 FreeSans 1120 90 0 0 la_oenb[125]
port 448 nsew signal input
flabel metal2 s 574976 -800 575088 480 0 FreeSans 1120 90 0 0 la_oenb[126]
port 449 nsew signal input
flabel metal2 s 578522 -800 578634 480 0 FreeSans 1120 90 0 0 la_oenb[127]
port 450 nsew signal input
flabel metal2 s 170732 -800 170844 480 0 FreeSans 1120 90 0 0 la_oenb[12]
port 451 nsew signal input
flabel metal2 s 174278 -800 174390 480 0 FreeSans 1120 90 0 0 la_oenb[13]
port 452 nsew signal input
flabel metal2 s 177824 -800 177936 480 0 FreeSans 1120 90 0 0 la_oenb[14]
port 453 nsew signal input
flabel metal2 s 181370 -800 181482 480 0 FreeSans 1120 90 0 0 la_oenb[15]
port 454 nsew signal input
flabel metal2 s 184916 -800 185028 480 0 FreeSans 1120 90 0 0 la_oenb[16]
port 455 nsew signal input
flabel metal2 s 188462 -800 188574 480 0 FreeSans 1120 90 0 0 la_oenb[17]
port 456 nsew signal input
flabel metal2 s 192008 -800 192120 480 0 FreeSans 1120 90 0 0 la_oenb[18]
port 457 nsew signal input
flabel metal2 s 195554 -800 195666 480 0 FreeSans 1120 90 0 0 la_oenb[19]
port 458 nsew signal input
flabel metal2 s 131726 -800 131838 480 0 FreeSans 1120 90 0 0 la_oenb[1]
port 459 nsew signal input
flabel metal2 s 199100 -800 199212 480 0 FreeSans 1120 90 0 0 la_oenb[20]
port 460 nsew signal input
flabel metal2 s 202646 -800 202758 480 0 FreeSans 1120 90 0 0 la_oenb[21]
port 461 nsew signal input
flabel metal2 s 206192 -800 206304 480 0 FreeSans 1120 90 0 0 la_oenb[22]
port 462 nsew signal input
flabel metal2 s 209738 -800 209850 480 0 FreeSans 1120 90 0 0 la_oenb[23]
port 463 nsew signal input
flabel metal2 s 213284 -800 213396 480 0 FreeSans 1120 90 0 0 la_oenb[24]
port 464 nsew signal input
flabel metal2 s 216830 -800 216942 480 0 FreeSans 1120 90 0 0 la_oenb[25]
port 465 nsew signal input
flabel metal2 s 220376 -800 220488 480 0 FreeSans 1120 90 0 0 la_oenb[26]
port 466 nsew signal input
flabel metal2 s 223922 -800 224034 480 0 FreeSans 1120 90 0 0 la_oenb[27]
port 467 nsew signal input
flabel metal2 s 227468 -800 227580 480 0 FreeSans 1120 90 0 0 la_oenb[28]
port 468 nsew signal input
flabel metal2 s 231014 -800 231126 480 0 FreeSans 1120 90 0 0 la_oenb[29]
port 469 nsew signal input
flabel metal2 s 135272 -800 135384 480 0 FreeSans 1120 90 0 0 la_oenb[2]
port 470 nsew signal input
flabel metal2 s 234560 -800 234672 480 0 FreeSans 1120 90 0 0 la_oenb[30]
port 471 nsew signal input
flabel metal2 s 238106 -800 238218 480 0 FreeSans 1120 90 0 0 la_oenb[31]
port 472 nsew signal input
flabel metal2 s 241652 -800 241764 480 0 FreeSans 1120 90 0 0 la_oenb[32]
port 473 nsew signal input
flabel metal2 s 245198 -800 245310 480 0 FreeSans 1120 90 0 0 la_oenb[33]
port 474 nsew signal input
flabel metal2 s 248744 -800 248856 480 0 FreeSans 1120 90 0 0 la_oenb[34]
port 475 nsew signal input
flabel metal2 s 252290 -800 252402 480 0 FreeSans 1120 90 0 0 la_oenb[35]
port 476 nsew signal input
flabel metal2 s 255836 -800 255948 480 0 FreeSans 1120 90 0 0 la_oenb[36]
port 477 nsew signal input
flabel metal2 s 259382 -800 259494 480 0 FreeSans 1120 90 0 0 la_oenb[37]
port 478 nsew signal input
flabel metal2 s 262928 -800 263040 480 0 FreeSans 1120 90 0 0 la_oenb[38]
port 479 nsew signal input
flabel metal2 s 266474 -800 266586 480 0 FreeSans 1120 90 0 0 la_oenb[39]
port 480 nsew signal input
flabel metal2 s 138818 -800 138930 480 0 FreeSans 1120 90 0 0 la_oenb[3]
port 481 nsew signal input
flabel metal2 s 270020 -800 270132 480 0 FreeSans 1120 90 0 0 la_oenb[40]
port 482 nsew signal input
flabel metal2 s 273566 -800 273678 480 0 FreeSans 1120 90 0 0 la_oenb[41]
port 483 nsew signal input
flabel metal2 s 277112 -800 277224 480 0 FreeSans 1120 90 0 0 la_oenb[42]
port 484 nsew signal input
flabel metal2 s 280658 -800 280770 480 0 FreeSans 1120 90 0 0 la_oenb[43]
port 485 nsew signal input
flabel metal2 s 284204 -800 284316 480 0 FreeSans 1120 90 0 0 la_oenb[44]
port 486 nsew signal input
flabel metal2 s 287750 -800 287862 480 0 FreeSans 1120 90 0 0 la_oenb[45]
port 487 nsew signal input
flabel metal2 s 291296 -800 291408 480 0 FreeSans 1120 90 0 0 la_oenb[46]
port 488 nsew signal input
flabel metal2 s 294842 -800 294954 480 0 FreeSans 1120 90 0 0 la_oenb[47]
port 489 nsew signal input
flabel metal2 s 298388 -800 298500 480 0 FreeSans 1120 90 0 0 la_oenb[48]
port 490 nsew signal input
flabel metal2 s 301934 -800 302046 480 0 FreeSans 1120 90 0 0 la_oenb[49]
port 491 nsew signal input
flabel metal2 s 142364 -800 142476 480 0 FreeSans 1120 90 0 0 la_oenb[4]
port 492 nsew signal input
flabel metal2 s 305480 -800 305592 480 0 FreeSans 1120 90 0 0 la_oenb[50]
port 493 nsew signal input
flabel metal2 s 309026 -800 309138 480 0 FreeSans 1120 90 0 0 la_oenb[51]
port 494 nsew signal input
flabel metal2 s 312572 -800 312684 480 0 FreeSans 1120 90 0 0 la_oenb[52]
port 495 nsew signal input
flabel metal2 s 316118 -800 316230 480 0 FreeSans 1120 90 0 0 la_oenb[53]
port 496 nsew signal input
flabel metal2 s 319664 -800 319776 480 0 FreeSans 1120 90 0 0 la_oenb[54]
port 497 nsew signal input
flabel metal2 s 323210 -800 323322 480 0 FreeSans 1120 90 0 0 la_oenb[55]
port 498 nsew signal input
flabel metal2 s 326756 -800 326868 480 0 FreeSans 1120 90 0 0 la_oenb[56]
port 499 nsew signal input
flabel metal2 s 330302 -800 330414 480 0 FreeSans 1120 90 0 0 la_oenb[57]
port 500 nsew signal input
flabel metal2 s 333848 -800 333960 480 0 FreeSans 1120 90 0 0 la_oenb[58]
port 501 nsew signal input
flabel metal2 s 337394 -800 337506 480 0 FreeSans 1120 90 0 0 la_oenb[59]
port 502 nsew signal input
flabel metal2 s 145910 -800 146022 480 0 FreeSans 1120 90 0 0 la_oenb[5]
port 503 nsew signal input
flabel metal2 s 340940 -800 341052 480 0 FreeSans 1120 90 0 0 la_oenb[60]
port 504 nsew signal input
flabel metal2 s 344486 -800 344598 480 0 FreeSans 1120 90 0 0 la_oenb[61]
port 505 nsew signal input
flabel metal2 s 348032 -800 348144 480 0 FreeSans 1120 90 0 0 la_oenb[62]
port 506 nsew signal input
flabel metal2 s 351578 -800 351690 480 0 FreeSans 1120 90 0 0 la_oenb[63]
port 507 nsew signal input
flabel metal2 s 355124 -800 355236 480 0 FreeSans 1120 90 0 0 la_oenb[64]
port 508 nsew signal input
flabel metal2 s 358670 -800 358782 480 0 FreeSans 1120 90 0 0 la_oenb[65]
port 509 nsew signal input
flabel metal2 s 362216 -800 362328 480 0 FreeSans 1120 90 0 0 la_oenb[66]
port 510 nsew signal input
flabel metal2 s 365762 -800 365874 480 0 FreeSans 1120 90 0 0 la_oenb[67]
port 511 nsew signal input
flabel metal2 s 369308 -800 369420 480 0 FreeSans 1120 90 0 0 la_oenb[68]
port 512 nsew signal input
flabel metal2 s 372854 -800 372966 480 0 FreeSans 1120 90 0 0 la_oenb[69]
port 513 nsew signal input
flabel metal2 s 149456 -800 149568 480 0 FreeSans 1120 90 0 0 la_oenb[6]
port 514 nsew signal input
flabel metal2 s 376400 -800 376512 480 0 FreeSans 1120 90 0 0 la_oenb[70]
port 515 nsew signal input
flabel metal2 s 379946 -800 380058 480 0 FreeSans 1120 90 0 0 la_oenb[71]
port 516 nsew signal input
flabel metal2 s 383492 -800 383604 480 0 FreeSans 1120 90 0 0 la_oenb[72]
port 517 nsew signal input
flabel metal2 s 387038 -800 387150 480 0 FreeSans 1120 90 0 0 la_oenb[73]
port 518 nsew signal input
flabel metal2 s 390584 -800 390696 480 0 FreeSans 1120 90 0 0 la_oenb[74]
port 519 nsew signal input
flabel metal2 s 394130 -800 394242 480 0 FreeSans 1120 90 0 0 la_oenb[75]
port 520 nsew signal input
flabel metal2 s 397676 -800 397788 480 0 FreeSans 1120 90 0 0 la_oenb[76]
port 521 nsew signal input
flabel metal2 s 401222 -800 401334 480 0 FreeSans 1120 90 0 0 la_oenb[77]
port 522 nsew signal input
flabel metal2 s 404768 -800 404880 480 0 FreeSans 1120 90 0 0 la_oenb[78]
port 523 nsew signal input
flabel metal2 s 408314 -800 408426 480 0 FreeSans 1120 90 0 0 la_oenb[79]
port 524 nsew signal input
flabel metal2 s 153002 -800 153114 480 0 FreeSans 1120 90 0 0 la_oenb[7]
port 525 nsew signal input
flabel metal2 s 411860 -800 411972 480 0 FreeSans 1120 90 0 0 la_oenb[80]
port 526 nsew signal input
flabel metal2 s 415406 -800 415518 480 0 FreeSans 1120 90 0 0 la_oenb[81]
port 527 nsew signal input
flabel metal2 s 418952 -800 419064 480 0 FreeSans 1120 90 0 0 la_oenb[82]
port 528 nsew signal input
flabel metal2 s 422498 -800 422610 480 0 FreeSans 1120 90 0 0 la_oenb[83]
port 529 nsew signal input
flabel metal2 s 426044 -800 426156 480 0 FreeSans 1120 90 0 0 la_oenb[84]
port 530 nsew signal input
flabel metal2 s 429590 -800 429702 480 0 FreeSans 1120 90 0 0 la_oenb[85]
port 531 nsew signal input
flabel metal2 s 433136 -800 433248 480 0 FreeSans 1120 90 0 0 la_oenb[86]
port 532 nsew signal input
flabel metal2 s 436682 -800 436794 480 0 FreeSans 1120 90 0 0 la_oenb[87]
port 533 nsew signal input
flabel metal2 s 440228 -800 440340 480 0 FreeSans 1120 90 0 0 la_oenb[88]
port 534 nsew signal input
flabel metal2 s 443774 -800 443886 480 0 FreeSans 1120 90 0 0 la_oenb[89]
port 535 nsew signal input
flabel metal2 s 156548 -800 156660 480 0 FreeSans 1120 90 0 0 la_oenb[8]
port 536 nsew signal input
flabel metal2 s 447320 -800 447432 480 0 FreeSans 1120 90 0 0 la_oenb[90]
port 537 nsew signal input
flabel metal2 s 450866 -800 450978 480 0 FreeSans 1120 90 0 0 la_oenb[91]
port 538 nsew signal input
flabel metal2 s 454412 -800 454524 480 0 FreeSans 1120 90 0 0 la_oenb[92]
port 539 nsew signal input
flabel metal2 s 457958 -800 458070 480 0 FreeSans 1120 90 0 0 la_oenb[93]
port 540 nsew signal input
flabel metal2 s 461504 -800 461616 480 0 FreeSans 1120 90 0 0 la_oenb[94]
port 541 nsew signal input
flabel metal2 s 465050 -800 465162 480 0 FreeSans 1120 90 0 0 la_oenb[95]
port 542 nsew signal input
flabel metal2 s 468596 -800 468708 480 0 FreeSans 1120 90 0 0 la_oenb[96]
port 543 nsew signal input
flabel metal2 s 472142 -800 472254 480 0 FreeSans 1120 90 0 0 la_oenb[97]
port 544 nsew signal input
flabel metal2 s 475688 -800 475800 480 0 FreeSans 1120 90 0 0 la_oenb[98]
port 545 nsew signal input
flabel metal2 s 479234 -800 479346 480 0 FreeSans 1120 90 0 0 la_oenb[99]
port 546 nsew signal input
flabel metal2 s 160094 -800 160206 480 0 FreeSans 1120 90 0 0 la_oenb[9]
port 547 nsew signal input
flabel metal2 s 579704 -800 579816 480 0 FreeSans 1120 90 0 0 user_clock2
port 548 nsew signal input
flabel metal2 s 580886 -800 580998 480 0 FreeSans 1120 90 0 0 user_irq[0]
port 549 nsew signal tristate
flabel metal2 s 582068 -800 582180 480 0 FreeSans 1120 90 0 0 user_irq[1]
port 550 nsew signal tristate
flabel metal2 s 583250 -800 583362 480 0 FreeSans 1120 90 0 0 user_irq[2]
port 551 nsew signal tristate
flabel metal3 s 582340 639784 584800 644584 0 FreeSans 1120 0 0 0 vccd1
port 552 nsew signal bidirectional
flabel metal3 s 582340 629784 584800 634584 0 FreeSans 1120 0 0 0 vccd1
port 553 nsew signal bidirectional
flabel metal3 s 0 643842 1660 648642 0 FreeSans 1120 0 0 0 vccd2
port 554 nsew signal bidirectional
flabel metal3 s 0 633842 1660 638642 0 FreeSans 1120 0 0 0 vccd2
port 555 nsew signal bidirectional
flabel metal3 s 582340 540562 584800 545362 0 FreeSans 1120 0 0 0 vdda1
port 556 nsew signal bidirectional
flabel metal3 s 582340 550562 584800 555362 0 FreeSans 1120 0 0 0 vdda1
port 557 nsew signal bidirectional
flabel metal3 s 582340 235230 584800 240030 0 FreeSans 1120 0 0 0 vdda1
port 558 nsew signal bidirectional
flabel metal3 s 582340 225230 584800 230030 0 FreeSans 1120 0 0 0 vdda1
port 559 nsew signal bidirectional
flabel metal3 s 0 204888 1660 209688 0 FreeSans 1120 0 0 0 vdda2
port 560 nsew signal bidirectional
flabel metal3 s 0 214888 1660 219688 0 FreeSans 1120 0 0 0 vdda2
port 561 nsew signal bidirectional
flabel metal3 s 520594 702340 525394 704800 0 FreeSans 1920 180 0 0 vssa1
port 562 nsew signal bidirectional
flabel metal3 s 510594 702340 515394 704800 0 FreeSans 1920 180 0 0 vssa1
port 563 nsew signal bidirectional
flabel metal3 s 582340 146830 584800 151630 0 FreeSans 1120 0 0 0 vssa1
port 564 nsew signal bidirectional
flabel metal3 s 582340 136830 584800 141630 0 FreeSans 1120 0 0 0 vssa1
port 565 nsew signal bidirectional
flabel metal3 s 0 559442 1660 564242 0 FreeSans 1120 0 0 0 vssa2
port 566 nsew signal bidirectional
flabel metal3 s 0 549442 1660 554242 0 FreeSans 1120 0 0 0 vssa2
port 567 nsew signal bidirectional
flabel metal3 s 582340 191430 584800 196230 0 FreeSans 1120 0 0 0 vssd1
port 568 nsew signal bidirectional
flabel metal3 s 582340 181430 584800 186230 0 FreeSans 1120 0 0 0 vssd1
port 569 nsew signal bidirectional
flabel metal3 s 0 172888 1660 177688 0 FreeSans 1120 0 0 0 vssd2
port 570 nsew signal bidirectional
flabel metal3 s 0 162888 1660 167688 0 FreeSans 1120 0 0 0 vssd2
port 571 nsew signal bidirectional
flabel metal2 s 524 -800 636 480 0 FreeSans 1120 90 0 0 wb_clk_i
port 572 nsew signal input
flabel metal2 s 1706 -800 1818 480 0 FreeSans 1120 90 0 0 wb_rst_i
port 573 nsew signal input
flabel metal2 s 2888 -800 3000 480 0 FreeSans 1120 90 0 0 wbs_ack_o
port 574 nsew signal tristate
flabel metal2 s 7616 -800 7728 480 0 FreeSans 1120 90 0 0 wbs_adr_i[0]
port 575 nsew signal input
flabel metal2 s 47804 -800 47916 480 0 FreeSans 1120 90 0 0 wbs_adr_i[10]
port 576 nsew signal input
flabel metal2 s 51350 -800 51462 480 0 FreeSans 1120 90 0 0 wbs_adr_i[11]
port 577 nsew signal input
flabel metal2 s 54896 -800 55008 480 0 FreeSans 1120 90 0 0 wbs_adr_i[12]
port 578 nsew signal input
flabel metal2 s 58442 -800 58554 480 0 FreeSans 1120 90 0 0 wbs_adr_i[13]
port 579 nsew signal input
flabel metal2 s 61988 -800 62100 480 0 FreeSans 1120 90 0 0 wbs_adr_i[14]
port 580 nsew signal input
flabel metal2 s 65534 -800 65646 480 0 FreeSans 1120 90 0 0 wbs_adr_i[15]
port 581 nsew signal input
flabel metal2 s 69080 -800 69192 480 0 FreeSans 1120 90 0 0 wbs_adr_i[16]
port 582 nsew signal input
flabel metal2 s 72626 -800 72738 480 0 FreeSans 1120 90 0 0 wbs_adr_i[17]
port 583 nsew signal input
flabel metal2 s 76172 -800 76284 480 0 FreeSans 1120 90 0 0 wbs_adr_i[18]
port 584 nsew signal input
flabel metal2 s 79718 -800 79830 480 0 FreeSans 1120 90 0 0 wbs_adr_i[19]
port 585 nsew signal input
flabel metal2 s 12344 -800 12456 480 0 FreeSans 1120 90 0 0 wbs_adr_i[1]
port 586 nsew signal input
flabel metal2 s 83264 -800 83376 480 0 FreeSans 1120 90 0 0 wbs_adr_i[20]
port 587 nsew signal input
flabel metal2 s 86810 -800 86922 480 0 FreeSans 1120 90 0 0 wbs_adr_i[21]
port 588 nsew signal input
flabel metal2 s 90356 -800 90468 480 0 FreeSans 1120 90 0 0 wbs_adr_i[22]
port 589 nsew signal input
flabel metal2 s 93902 -800 94014 480 0 FreeSans 1120 90 0 0 wbs_adr_i[23]
port 590 nsew signal input
flabel metal2 s 97448 -800 97560 480 0 FreeSans 1120 90 0 0 wbs_adr_i[24]
port 591 nsew signal input
flabel metal2 s 100994 -800 101106 480 0 FreeSans 1120 90 0 0 wbs_adr_i[25]
port 592 nsew signal input
flabel metal2 s 104540 -800 104652 480 0 FreeSans 1120 90 0 0 wbs_adr_i[26]
port 593 nsew signal input
flabel metal2 s 108086 -800 108198 480 0 FreeSans 1120 90 0 0 wbs_adr_i[27]
port 594 nsew signal input
flabel metal2 s 111632 -800 111744 480 0 FreeSans 1120 90 0 0 wbs_adr_i[28]
port 595 nsew signal input
flabel metal2 s 115178 -800 115290 480 0 FreeSans 1120 90 0 0 wbs_adr_i[29]
port 596 nsew signal input
flabel metal2 s 17072 -800 17184 480 0 FreeSans 1120 90 0 0 wbs_adr_i[2]
port 597 nsew signal input
flabel metal2 s 118724 -800 118836 480 0 FreeSans 1120 90 0 0 wbs_adr_i[30]
port 598 nsew signal input
flabel metal2 s 122270 -800 122382 480 0 FreeSans 1120 90 0 0 wbs_adr_i[31]
port 599 nsew signal input
flabel metal2 s 21800 -800 21912 480 0 FreeSans 1120 90 0 0 wbs_adr_i[3]
port 600 nsew signal input
flabel metal2 s 26528 -800 26640 480 0 FreeSans 1120 90 0 0 wbs_adr_i[4]
port 601 nsew signal input
flabel metal2 s 30074 -800 30186 480 0 FreeSans 1120 90 0 0 wbs_adr_i[5]
port 602 nsew signal input
flabel metal2 s 33620 -800 33732 480 0 FreeSans 1120 90 0 0 wbs_adr_i[6]
port 603 nsew signal input
flabel metal2 s 37166 -800 37278 480 0 FreeSans 1120 90 0 0 wbs_adr_i[7]
port 604 nsew signal input
flabel metal2 s 40712 -800 40824 480 0 FreeSans 1120 90 0 0 wbs_adr_i[8]
port 605 nsew signal input
flabel metal2 s 44258 -800 44370 480 0 FreeSans 1120 90 0 0 wbs_adr_i[9]
port 606 nsew signal input
flabel metal2 s 4070 -800 4182 480 0 FreeSans 1120 90 0 0 wbs_cyc_i
port 607 nsew signal input
flabel metal2 s 8798 -800 8910 480 0 FreeSans 1120 90 0 0 wbs_dat_i[0]
port 608 nsew signal input
flabel metal2 s 48986 -800 49098 480 0 FreeSans 1120 90 0 0 wbs_dat_i[10]
port 609 nsew signal input
flabel metal2 s 52532 -800 52644 480 0 FreeSans 1120 90 0 0 wbs_dat_i[11]
port 610 nsew signal input
flabel metal2 s 56078 -800 56190 480 0 FreeSans 1120 90 0 0 wbs_dat_i[12]
port 611 nsew signal input
flabel metal2 s 59624 -800 59736 480 0 FreeSans 1120 90 0 0 wbs_dat_i[13]
port 612 nsew signal input
flabel metal2 s 63170 -800 63282 480 0 FreeSans 1120 90 0 0 wbs_dat_i[14]
port 613 nsew signal input
flabel metal2 s 66716 -800 66828 480 0 FreeSans 1120 90 0 0 wbs_dat_i[15]
port 614 nsew signal input
flabel metal2 s 70262 -800 70374 480 0 FreeSans 1120 90 0 0 wbs_dat_i[16]
port 615 nsew signal input
flabel metal2 s 73808 -800 73920 480 0 FreeSans 1120 90 0 0 wbs_dat_i[17]
port 616 nsew signal input
flabel metal2 s 77354 -800 77466 480 0 FreeSans 1120 90 0 0 wbs_dat_i[18]
port 617 nsew signal input
flabel metal2 s 80900 -800 81012 480 0 FreeSans 1120 90 0 0 wbs_dat_i[19]
port 618 nsew signal input
flabel metal2 s 13526 -800 13638 480 0 FreeSans 1120 90 0 0 wbs_dat_i[1]
port 619 nsew signal input
flabel metal2 s 84446 -800 84558 480 0 FreeSans 1120 90 0 0 wbs_dat_i[20]
port 620 nsew signal input
flabel metal2 s 87992 -800 88104 480 0 FreeSans 1120 90 0 0 wbs_dat_i[21]
port 621 nsew signal input
flabel metal2 s 91538 -800 91650 480 0 FreeSans 1120 90 0 0 wbs_dat_i[22]
port 622 nsew signal input
flabel metal2 s 95084 -800 95196 480 0 FreeSans 1120 90 0 0 wbs_dat_i[23]
port 623 nsew signal input
flabel metal2 s 98630 -800 98742 480 0 FreeSans 1120 90 0 0 wbs_dat_i[24]
port 624 nsew signal input
flabel metal2 s 102176 -800 102288 480 0 FreeSans 1120 90 0 0 wbs_dat_i[25]
port 625 nsew signal input
flabel metal2 s 105722 -800 105834 480 0 FreeSans 1120 90 0 0 wbs_dat_i[26]
port 626 nsew signal input
flabel metal2 s 109268 -800 109380 480 0 FreeSans 1120 90 0 0 wbs_dat_i[27]
port 627 nsew signal input
flabel metal2 s 112814 -800 112926 480 0 FreeSans 1120 90 0 0 wbs_dat_i[28]
port 628 nsew signal input
flabel metal2 s 116360 -800 116472 480 0 FreeSans 1120 90 0 0 wbs_dat_i[29]
port 629 nsew signal input
flabel metal2 s 18254 -800 18366 480 0 FreeSans 1120 90 0 0 wbs_dat_i[2]
port 630 nsew signal input
flabel metal2 s 119906 -800 120018 480 0 FreeSans 1120 90 0 0 wbs_dat_i[30]
port 631 nsew signal input
flabel metal2 s 123452 -800 123564 480 0 FreeSans 1120 90 0 0 wbs_dat_i[31]
port 632 nsew signal input
flabel metal2 s 22982 -800 23094 480 0 FreeSans 1120 90 0 0 wbs_dat_i[3]
port 633 nsew signal input
flabel metal2 s 27710 -800 27822 480 0 FreeSans 1120 90 0 0 wbs_dat_i[4]
port 634 nsew signal input
flabel metal2 s 31256 -800 31368 480 0 FreeSans 1120 90 0 0 wbs_dat_i[5]
port 635 nsew signal input
flabel metal2 s 34802 -800 34914 480 0 FreeSans 1120 90 0 0 wbs_dat_i[6]
port 636 nsew signal input
flabel metal2 s 38348 -800 38460 480 0 FreeSans 1120 90 0 0 wbs_dat_i[7]
port 637 nsew signal input
flabel metal2 s 41894 -800 42006 480 0 FreeSans 1120 90 0 0 wbs_dat_i[8]
port 638 nsew signal input
flabel metal2 s 45440 -800 45552 480 0 FreeSans 1120 90 0 0 wbs_dat_i[9]
port 639 nsew signal input
flabel metal2 s 9980 -800 10092 480 0 FreeSans 1120 90 0 0 wbs_dat_o[0]
port 640 nsew signal tristate
flabel metal2 s 50168 -800 50280 480 0 FreeSans 1120 90 0 0 wbs_dat_o[10]
port 641 nsew signal tristate
flabel metal2 s 53714 -800 53826 480 0 FreeSans 1120 90 0 0 wbs_dat_o[11]
port 642 nsew signal tristate
flabel metal2 s 57260 -800 57372 480 0 FreeSans 1120 90 0 0 wbs_dat_o[12]
port 643 nsew signal tristate
flabel metal2 s 60806 -800 60918 480 0 FreeSans 1120 90 0 0 wbs_dat_o[13]
port 644 nsew signal tristate
flabel metal2 s 64352 -800 64464 480 0 FreeSans 1120 90 0 0 wbs_dat_o[14]
port 645 nsew signal tristate
flabel metal2 s 67898 -800 68010 480 0 FreeSans 1120 90 0 0 wbs_dat_o[15]
port 646 nsew signal tristate
flabel metal2 s 71444 -800 71556 480 0 FreeSans 1120 90 0 0 wbs_dat_o[16]
port 647 nsew signal tristate
flabel metal2 s 74990 -800 75102 480 0 FreeSans 1120 90 0 0 wbs_dat_o[17]
port 648 nsew signal tristate
flabel metal2 s 78536 -800 78648 480 0 FreeSans 1120 90 0 0 wbs_dat_o[18]
port 649 nsew signal tristate
flabel metal2 s 82082 -800 82194 480 0 FreeSans 1120 90 0 0 wbs_dat_o[19]
port 650 nsew signal tristate
flabel metal2 s 14708 -800 14820 480 0 FreeSans 1120 90 0 0 wbs_dat_o[1]
port 651 nsew signal tristate
flabel metal2 s 85628 -800 85740 480 0 FreeSans 1120 90 0 0 wbs_dat_o[20]
port 652 nsew signal tristate
flabel metal2 s 89174 -800 89286 480 0 FreeSans 1120 90 0 0 wbs_dat_o[21]
port 653 nsew signal tristate
flabel metal2 s 92720 -800 92832 480 0 FreeSans 1120 90 0 0 wbs_dat_o[22]
port 654 nsew signal tristate
flabel metal2 s 96266 -800 96378 480 0 FreeSans 1120 90 0 0 wbs_dat_o[23]
port 655 nsew signal tristate
flabel metal2 s 99812 -800 99924 480 0 FreeSans 1120 90 0 0 wbs_dat_o[24]
port 656 nsew signal tristate
flabel metal2 s 103358 -800 103470 480 0 FreeSans 1120 90 0 0 wbs_dat_o[25]
port 657 nsew signal tristate
flabel metal2 s 106904 -800 107016 480 0 FreeSans 1120 90 0 0 wbs_dat_o[26]
port 658 nsew signal tristate
flabel metal2 s 110450 -800 110562 480 0 FreeSans 1120 90 0 0 wbs_dat_o[27]
port 659 nsew signal tristate
flabel metal2 s 113996 -800 114108 480 0 FreeSans 1120 90 0 0 wbs_dat_o[28]
port 660 nsew signal tristate
flabel metal2 s 117542 -800 117654 480 0 FreeSans 1120 90 0 0 wbs_dat_o[29]
port 661 nsew signal tristate
flabel metal2 s 19436 -800 19548 480 0 FreeSans 1120 90 0 0 wbs_dat_o[2]
port 662 nsew signal tristate
flabel metal2 s 121088 -800 121200 480 0 FreeSans 1120 90 0 0 wbs_dat_o[30]
port 663 nsew signal tristate
flabel metal2 s 124634 -800 124746 480 0 FreeSans 1120 90 0 0 wbs_dat_o[31]
port 664 nsew signal tristate
flabel metal2 s 24164 -800 24276 480 0 FreeSans 1120 90 0 0 wbs_dat_o[3]
port 665 nsew signal tristate
flabel metal2 s 28892 -800 29004 480 0 FreeSans 1120 90 0 0 wbs_dat_o[4]
port 666 nsew signal tristate
flabel metal2 s 32438 -800 32550 480 0 FreeSans 1120 90 0 0 wbs_dat_o[5]
port 667 nsew signal tristate
flabel metal2 s 35984 -800 36096 480 0 FreeSans 1120 90 0 0 wbs_dat_o[6]
port 668 nsew signal tristate
flabel metal2 s 39530 -800 39642 480 0 FreeSans 1120 90 0 0 wbs_dat_o[7]
port 669 nsew signal tristate
flabel metal2 s 43076 -800 43188 480 0 FreeSans 1120 90 0 0 wbs_dat_o[8]
port 670 nsew signal tristate
flabel metal2 s 46622 -800 46734 480 0 FreeSans 1120 90 0 0 wbs_dat_o[9]
port 671 nsew signal tristate
flabel metal2 s 11162 -800 11274 480 0 FreeSans 1120 90 0 0 wbs_sel_i[0]
port 672 nsew signal input
flabel metal2 s 15890 -800 16002 480 0 FreeSans 1120 90 0 0 wbs_sel_i[1]
port 673 nsew signal input
flabel metal2 s 20618 -800 20730 480 0 FreeSans 1120 90 0 0 wbs_sel_i[2]
port 674 nsew signal input
flabel metal2 s 25346 -800 25458 480 0 FreeSans 1120 90 0 0 wbs_sel_i[3]
port 675 nsew signal input
flabel metal2 s 5252 -800 5364 480 0 FreeSans 1120 90 0 0 wbs_stb_i
port 676 nsew signal input
flabel metal2 s 6434 -800 6546 480 0 FreeSans 1120 90 0 0 wbs_we_i
port 677 nsew signal input
flabel metal1 509928 469744 510126 470206 3 FreeSans 1600 0 0 0 bandgaptop_flat_io_0/bandgaptop_flat_0/porst
flabel metal1 514250 449142 514926 453810 3 FreeSans 1600 0 0 0 bandgaptop_flat_io_0/bandgaptop_flat_0/Vbg
flabel metal2 506154 470482 506224 472264 3 FreeSans 800 0 0 0 bandgaptop_flat_io_0/bandgaptop_flat_0/ampcurrentsource_0/Vq
flabel metal2 506364 470482 506434 472264 3 FreeSans 800 0 0 0 bandgaptop_flat_io_0/bandgaptop_flat_0/ampcurrentsource_0/Vx
flabel locali 507124 471322 507152 471404 3 FreeSans 800 0 0 0 bandgaptop_flat_io_0/bandgaptop_flat_0/ampcurrentsource_0/GND!
flabel metal2 502864 465496 502988 465512 7 FreeSans 800 0 0 0 bandgaptop_flat_io_0/bandgaptop_flat_0/amplifier_0/VDD!
flabel metal2 506092 464842 506216 464858 7 FreeSans 800 0 0 0 bandgaptop_flat_io_0/bandgaptop_flat_0/amplifier_0/Vq
flabel metal2 508352 464900 508432 464916 7 FreeSans 800 0 0 0 bandgaptop_flat_io_0/bandgaptop_flat_0/amplifier_0/Va
flabel metal2 508212 465672 508292 465688 7 FreeSans 800 0 0 0 bandgaptop_flat_io_0/bandgaptop_flat_0/amplifier_0/Vb
flabel metal2 505796 464088 506062 464182 7 FreeSans 800 0 0 0 bandgaptop_flat_io_0/bandgaptop_flat_0/amplifier_0/Vgate
flabel metal2 505796 465812 506062 465906 7 FreeSans 800 0 0 0 bandgaptop_flat_io_0/bandgaptop_flat_0/amplifier_0/Vgate
flabel metal1 505810 467230 505902 467264 7 FreeSans 800 0 0 0 bandgaptop_flat_io_0/bandgaptop_flat_0/amplifier_0/vg
flabel metal2 502664 463142 502788 463164 7 FreeSans 800 0 0 0 bandgaptop_flat_io_0/bandgaptop_flat_0/amplifier_0/Vx
flabel psubdiffcont 506468 468286 508068 468386 7 FreeSans 800 0 0 0 bandgaptop_flat_io_0/bandgaptop_flat_0/amplifier_0/GND!
flabel psubdiff 508068 462736 508168 462936 7 FreeSans 800 180 0 0 bandgaptop_flat_io_0/bandgaptop_flat_0/amplifier_0/GND!
rlabel via1 502844 459024 502888 459070 7 bandgaptop_flat_io_0/bandgaptop_flat_0/currentmirror_0/Vgate
rlabel metal3 502488 458214 502606 458348 7 bandgaptop_flat_io_0/bandgaptop_flat_0/currentmirror_0/VDD!
flabel metal1 511028 451242 511128 451542 7 FreeSans 1600 0 0 0 bandgaptop_flat_io_0/bandgaptop_flat_0/currentmirror_0/Vbg
flabel metal2 511628 451342 511728 451542 7 FreeSans 1600 0 0 0 bandgaptop_flat_io_0/bandgaptop_flat_0/currentmirror_0/Vb
flabel via2 512228 451342 512328 451542 7 FreeSans 1600 0 0 0 bandgaptop_flat_io_0/bandgaptop_flat_0/currentmirror_0/Va
flabel metal2 522926 449498 523358 450068 3 FreeSans 800 90 0 0 bandgaptop_flat_io_0/bandgaptop_flat_0/bandgapcorev3_0/VbEnd
flabel metal2 516190 448680 516622 449250 3 FreeSans 800 90 0 0 bandgaptop_flat_io_0/bandgaptop_flat_0/bandgapcorev3_0/VbgEnd
flabel metal2 522126 450316 523358 450886 3 FreeSans 800 90 0 0 bandgaptop_flat_io_0/bandgaptop_flat_0/bandgapcorev3_0/VaEnd
flabel metal2 515924 440450 516616 441142 3 FreeSans 1600 90 0 0 bandgaptop_flat_io_0/bandgaptop_flat_0/bandgapcorev3_0/Vbg
flabel metal2 515918 438808 516622 439512 3 FreeSans 1600 90 0 0 bandgaptop_flat_io_0/bandgaptop_flat_0/bandgapcorev3_0/Vb
flabel metal1 515352 439626 515924 440330 5 FreeSans 1600 0 0 0 bandgaptop_flat_io_0/bandgaptop_flat_0/bandgapcorev3_0/Va
rlabel psubdiffcont 500368 432068 501368 475308 3 bandgaptop_flat_io_0/bandgaptop_flat_0/GND
rlabel metal3 502426 470508 502848 471218 3 bandgaptop_flat_io_0/bandgaptop_flat_0/VDD
flabel metal2 503646 438210 504594 439346 1 FreeSans 1600 0 0 0 bandgaptop_flat_io_0/bandgaptop_flat_0/bandgapcorev3_0/Vbneg
flabel locali 503970 437706 504074 437954 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[0,0]/Emitter
flabel locali 504596 437794 504645 437895 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[0,0]/Collector
flabel locali 504446 437800 504486 437918 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[0,0]/Base
flabel locali 503970 436418 504074 436666 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[0,1]/Emitter
flabel locali 504596 436506 504645 436607 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[0,1]/Collector
flabel locali 504446 436512 504486 436630 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[0,1]/Base
flabel locali 503970 435130 504074 435378 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[0,2]/Emitter
flabel locali 504596 435218 504645 435319 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[0,2]/Collector
flabel locali 504446 435224 504486 435342 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[0,2]/Base
flabel locali 503970 433842 504074 434090 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[0,3]/Emitter
flabel locali 504596 433930 504645 434031 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[0,3]/Collector
flabel locali 504446 433936 504486 434054 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[0,3]/Base
flabel locali 503970 432554 504074 432802 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[0,4]/Emitter
flabel locali 504596 432642 504645 432743 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[0,4]/Collector
flabel locali 504446 432648 504486 432766 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[0,4]/Base
flabel locali 505258 437706 505362 437954 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[1,0]/Emitter
flabel locali 505884 437794 505933 437895 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[1,0]/Collector
flabel locali 505734 437800 505774 437918 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[1,0]/Base
flabel locali 505258 436418 505362 436666 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[1,1]/Emitter
flabel locali 505884 436506 505933 436607 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[1,1]/Collector
flabel locali 505734 436512 505774 436630 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[1,1]/Base
flabel locali 505258 435130 505362 435378 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[1,2]/Emitter
flabel locali 505884 435218 505933 435319 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[1,2]/Collector
flabel locali 505734 435224 505774 435342 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[1,2]/Base
flabel locali 505258 433842 505362 434090 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[1,3]/Emitter
flabel locali 505884 433930 505933 434031 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[1,3]/Collector
flabel locali 505734 433936 505774 434054 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[1,3]/Base
flabel locali 505258 432554 505362 432802 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[1,4]/Emitter
flabel locali 505884 432642 505933 432743 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[1,4]/Collector
flabel locali 505734 432648 505774 432766 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[1,4]/Base
flabel locali 506546 437706 506650 437954 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[2,0]/Emitter
flabel locali 507172 437794 507221 437895 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[2,0]/Collector
flabel locali 507022 437800 507062 437918 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[2,0]/Base
flabel locali 506546 436418 506650 436666 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[2,1]/Emitter
flabel locali 507172 436506 507221 436607 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[2,1]/Collector
flabel locali 507022 436512 507062 436630 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[2,1]/Base
flabel locali 506546 435130 506650 435378 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[2,2]/Emitter
flabel locali 507172 435218 507221 435319 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[2,2]/Collector
flabel locali 507022 435224 507062 435342 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[2,2]/Base
flabel locali 506546 433842 506650 434090 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[2,3]/Emitter
flabel locali 507172 433930 507221 434031 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[2,3]/Collector
flabel locali 507022 433936 507062 434054 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[2,3]/Base
flabel locali 506546 432554 506650 432802 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[2,4]/Emitter
flabel locali 507172 432642 507221 432743 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[2,4]/Collector
flabel locali 507022 432648 507062 432766 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[2,4]/Base
flabel locali 507834 437706 507938 437954 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[3,0]/Emitter
flabel locali 508460 437794 508509 437895 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[3,0]/Collector
flabel locali 508310 437800 508350 437918 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[3,0]/Base
flabel locali 507834 436418 507938 436666 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[3,1]/Emitter
flabel locali 508460 436506 508509 436607 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[3,1]/Collector
flabel locali 508310 436512 508350 436630 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[3,1]/Base
flabel locali 507834 435130 507938 435378 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[3,2]/Emitter
flabel locali 508460 435218 508509 435319 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[3,2]/Collector
flabel locali 508310 435224 508350 435342 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[3,2]/Base
flabel locali 507834 433842 507938 434090 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[3,3]/Emitter
flabel locali 508460 433930 508509 434031 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[3,3]/Collector
flabel locali 508310 433936 508350 434054 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[3,3]/Base
flabel locali 507834 432554 507938 432802 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[3,4]/Emitter
flabel locali 508460 432642 508509 432743 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[3,4]/Collector
flabel locali 508310 432648 508350 432766 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[3,4]/Base
flabel locali 509122 437706 509226 437954 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4,0]/Emitter
flabel locali 509748 437794 509797 437895 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4,0]/Collector
flabel locali 509598 437800 509638 437918 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4,0]/Base
flabel locali 509122 436418 509226 436666 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4,1]/Emitter
flabel locali 509748 436506 509797 436607 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4,1]/Collector
flabel locali 509598 436512 509638 436630 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4,1]/Base
flabel locali 509122 435130 509226 435378 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4,2]/Emitter
flabel locali 509748 435218 509797 435319 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4,2]/Collector
flabel locali 509598 435224 509638 435342 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4,2]/Base
flabel locali 509122 433842 509226 434090 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4,3]/Emitter
flabel locali 509748 433930 509797 434031 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4,3]/Collector
flabel locali 509598 433936 509638 434054 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4,3]/Base
flabel locali 509122 432554 509226 432802 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4,4]/Emitter
flabel locali 509748 432642 509797 432743 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4,4]/Collector
flabel locali 509598 432648 509638 432766 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[4,4]/Base
flabel locali 510410 437706 510514 437954 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[5,0]/Emitter
flabel locali 511036 437794 511085 437895 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[5,0]/Collector
flabel locali 510886 437800 510926 437918 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[5,0]/Base
flabel locali 510410 436418 510514 436666 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[5,1]/Emitter
flabel locali 511036 436506 511085 436607 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[5,1]/Collector
flabel locali 510886 436512 510926 436630 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[5,1]/Base
flabel locali 510410 435130 510514 435378 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[5,2]/Emitter
flabel locali 511036 435218 511085 435319 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[5,2]/Collector
flabel locali 510886 435224 510926 435342 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[5,2]/Base
flabel locali 510410 433842 510514 434090 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[5,3]/Emitter
flabel locali 511036 433930 511085 434031 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[5,3]/Collector
flabel locali 510886 433936 510926 434054 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[5,3]/Base
flabel locali 510410 432554 510514 432802 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[5,4]/Emitter
flabel locali 511036 432642 511085 432743 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[5,4]/Collector
flabel locali 510886 432648 510926 432766 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[5,4]/Base
flabel locali 511698 437706 511802 437954 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[6,0]/Emitter
flabel locali 512324 437794 512373 437895 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[6,0]/Collector
flabel locali 512174 437800 512214 437918 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[6,0]/Base
flabel locali 511698 436418 511802 436666 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[6,1]/Emitter
flabel locali 512324 436506 512373 436607 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[6,1]/Collector
flabel locali 512174 436512 512214 436630 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[6,1]/Base
flabel locali 511698 435130 511802 435378 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[6,2]/Emitter
flabel locali 512324 435218 512373 435319 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[6,2]/Collector
flabel locali 512174 435224 512214 435342 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[6,2]/Base
flabel locali 511698 433842 511802 434090 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[6,3]/Emitter
flabel locali 512324 433930 512373 434031 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[6,3]/Collector
flabel locali 512174 433936 512214 434054 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[6,3]/Base
flabel locali 511698 432554 511802 432802 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[6,4]/Emitter
flabel locali 512324 432642 512373 432743 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[6,4]/Collector
flabel locali 512174 432648 512214 432766 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[6,4]/Base
flabel locali 512986 437706 513090 437954 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[7,0]/Emitter
flabel locali 513612 437794 513661 437895 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[7,0]/Collector
flabel locali 513462 437800 513502 437918 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[7,0]/Base
flabel locali 512986 436418 513090 436666 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[7,1]/Emitter
flabel locali 513612 436506 513661 436607 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[7,1]/Collector
flabel locali 513462 436512 513502 436630 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[7,1]/Base
flabel locali 512986 435130 513090 435378 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[7,2]/Emitter
flabel locali 513612 435218 513661 435319 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[7,2]/Collector
flabel locali 513462 435224 513502 435342 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[7,2]/Base
flabel locali 512986 433842 513090 434090 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[7,3]/Emitter
flabel locali 513612 433930 513661 434031 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[7,3]/Collector
flabel locali 513462 433936 513502 434054 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[7,3]/Base
flabel locali 512986 432554 513090 432802 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[7,4]/Emitter
flabel locali 513612 432642 513661 432743 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[7,4]/Collector
flabel locali 513462 432648 513502 432766 0 FreeSans 400 0 0 0 bandgaptop_flat_io_0/sky130_fd_pr__rf_pnp_05v5_W3p40L3p40_0[7,4]/Base
<< end >>
