magic
tech sky130A
magscale 1 2
timestamp 1622327848
<< locali >>
rect 562528 494355 562562 494414
rect 563044 494355 563078 494414
rect 563560 494355 563594 494414
rect 564076 494355 564110 494414
rect 564592 494355 564626 494414
rect 565108 494355 565142 494414
rect 565624 494355 565658 494414
rect 566140 494355 566174 494414
rect 566656 494355 566690 494414
rect 567172 494355 567206 494414
rect 572688 494398 572722 494448
rect 573204 494398 573238 494448
rect 573720 494398 573754 494448
rect 574236 494398 574270 494448
rect 574752 494398 574786 494448
rect 575268 494398 575302 494448
rect 575784 494398 575818 494448
rect 576300 494398 576334 494448
rect 576816 494398 576850 494448
rect 577332 494398 577366 494448
rect 572429 494364 572476 494398
rect 572660 494364 577626 494398
rect 562270 494321 567234 494355
rect 567418 494321 567464 494355
rect 562528 454053 562562 454112
rect 563044 454053 563078 454112
rect 563560 454053 563594 454112
rect 564076 454053 564110 454112
rect 564592 454053 564626 454112
rect 565108 454053 565142 454112
rect 565624 454053 565658 454112
rect 566140 454053 566174 454112
rect 566656 454053 566690 454112
rect 567172 454053 567206 454112
rect 572688 454096 572722 454146
rect 573204 454096 573238 454146
rect 573720 454096 573754 454146
rect 574236 454096 574270 454146
rect 574752 454096 574786 454146
rect 575268 454096 575302 454146
rect 575784 454096 575818 454146
rect 576300 454096 576334 454146
rect 576816 454096 576850 454146
rect 577332 454096 577366 454146
rect 572429 454062 572476 454096
rect 572660 454062 577626 454096
rect 562270 454019 567234 454053
rect 567418 454019 567464 454053
<< metal1 >>
rect 562150 495742 567584 495775
rect 562150 495662 562480 495742
rect 562560 495662 562640 495742
rect 562720 495662 562800 495742
rect 562880 495662 562960 495742
rect 563040 495662 563120 495742
rect 563200 495662 563280 495742
rect 563360 495662 563440 495742
rect 563520 495662 563600 495742
rect 563680 495662 563760 495742
rect 563840 495662 563920 495742
rect 564000 495662 564080 495742
rect 564160 495662 564240 495742
rect 564320 495662 564400 495742
rect 564480 495662 564560 495742
rect 564640 495662 564720 495742
rect 564800 495662 564880 495742
rect 564960 495662 565040 495742
rect 565120 495662 565200 495742
rect 565280 495662 565360 495742
rect 565440 495662 565520 495742
rect 565600 495662 565680 495742
rect 565760 495662 565840 495742
rect 565920 495662 566000 495742
rect 566080 495662 566160 495742
rect 566240 495662 566320 495742
rect 566400 495662 566480 495742
rect 566560 495662 566640 495742
rect 566720 495662 566800 495742
rect 566880 495662 566960 495742
rect 567040 495662 567120 495742
rect 567200 495662 567280 495742
rect 567360 495662 567584 495742
rect 562150 495582 567584 495662
rect 562150 495502 562480 495582
rect 562560 495502 562640 495582
rect 562720 495502 562800 495582
rect 562880 495502 562960 495582
rect 563040 495502 563120 495582
rect 563200 495502 563280 495582
rect 563360 495502 563440 495582
rect 563520 495502 563600 495582
rect 563680 495502 563760 495582
rect 563840 495502 563920 495582
rect 564000 495502 564080 495582
rect 564160 495502 564240 495582
rect 564320 495502 564400 495582
rect 564480 495502 564560 495582
rect 564640 495502 564720 495582
rect 564800 495502 564880 495582
rect 564960 495502 565040 495582
rect 565120 495502 565200 495582
rect 565280 495502 565360 495582
rect 565440 495502 565520 495582
rect 565600 495502 565680 495582
rect 565760 495502 565840 495582
rect 565920 495502 566000 495582
rect 566080 495502 566160 495582
rect 566240 495502 566320 495582
rect 566400 495502 566480 495582
rect 566560 495502 566640 495582
rect 566720 495502 566800 495582
rect 566880 495502 566960 495582
rect 567040 495502 567120 495582
rect 567200 495502 567280 495582
rect 567360 495502 567584 495582
rect 562150 495474 567584 495502
rect 562150 494363 562196 495474
rect 562522 495402 562568 495474
rect 563038 495402 563084 495474
rect 563554 495402 563600 495474
rect 564070 495402 564116 495474
rect 564586 495402 564632 495474
rect 565102 495402 565148 495474
rect 565618 495402 565664 495474
rect 566134 495402 566180 495474
rect 566650 495402 566696 495474
rect 567166 495402 567212 495474
rect 562264 494277 562310 495402
rect 562780 494277 562826 495402
rect 563296 494277 563342 495402
rect 563812 494277 563858 495402
rect 564328 494277 564374 495402
rect 564844 494277 564890 495402
rect 565360 494277 565406 495402
rect 565876 494277 565922 495402
rect 566392 494277 566438 495402
rect 566908 494277 566954 495402
rect 567424 494277 567470 495402
rect 567538 494375 567584 495474
rect 572310 495742 577744 495775
rect 572310 495662 572640 495742
rect 572720 495662 572800 495742
rect 572880 495662 572960 495742
rect 573040 495662 573120 495742
rect 573200 495662 573280 495742
rect 573360 495662 573440 495742
rect 573520 495662 573600 495742
rect 573680 495662 573760 495742
rect 573840 495662 573920 495742
rect 574000 495662 574080 495742
rect 574160 495662 574240 495742
rect 574320 495662 574400 495742
rect 574480 495662 574560 495742
rect 574640 495662 574720 495742
rect 574800 495662 574880 495742
rect 574960 495662 575040 495742
rect 575120 495662 575200 495742
rect 575280 495662 575360 495742
rect 575440 495662 575520 495742
rect 575600 495662 575680 495742
rect 575760 495662 575840 495742
rect 575920 495662 576000 495742
rect 576080 495662 576160 495742
rect 576240 495662 576320 495742
rect 576400 495662 576480 495742
rect 576560 495662 576640 495742
rect 576720 495662 576800 495742
rect 576880 495662 576960 495742
rect 577040 495662 577120 495742
rect 577200 495662 577280 495742
rect 577360 495662 577440 495742
rect 577520 495662 577744 495742
rect 572310 495582 577744 495662
rect 572310 495502 572640 495582
rect 572720 495502 572800 495582
rect 572880 495502 572960 495582
rect 573040 495502 573120 495582
rect 573200 495502 573280 495582
rect 573360 495502 573440 495582
rect 573520 495502 573600 495582
rect 573680 495502 573760 495582
rect 573840 495502 573920 495582
rect 574000 495502 574080 495582
rect 574160 495502 574240 495582
rect 574320 495502 574400 495582
rect 574480 495502 574560 495582
rect 574640 495502 574720 495582
rect 574800 495502 574880 495582
rect 574960 495502 575040 495582
rect 575120 495502 575200 495582
rect 575280 495502 575360 495582
rect 575440 495502 575520 495582
rect 575600 495502 575680 495582
rect 575760 495502 575840 495582
rect 575920 495502 576000 495582
rect 576080 495502 576160 495582
rect 576240 495502 576320 495582
rect 576400 495502 576480 495582
rect 576560 495502 576640 495582
rect 576720 495502 576800 495582
rect 576880 495502 576960 495582
rect 577040 495502 577120 495582
rect 577200 495502 577280 495582
rect 577360 495502 577440 495582
rect 577520 495502 577744 495582
rect 572310 495474 577744 495502
rect 572310 495392 572356 495474
rect 572424 494292 572470 495436
rect 572688 495424 572722 495474
rect 572940 494292 572986 495436
rect 573204 495424 573238 495474
rect 573456 494292 573502 495436
rect 573720 495424 573754 495474
rect 573972 494292 574018 495436
rect 574236 495424 574270 495474
rect 574488 494292 574534 495436
rect 574752 495424 574786 495474
rect 575004 494292 575050 495436
rect 575268 495424 575302 495474
rect 575520 494292 575566 495436
rect 575784 495424 575818 495474
rect 576036 494292 576082 495436
rect 576300 495424 576334 495474
rect 576552 494292 576598 495436
rect 576816 495424 576850 495474
rect 577068 494292 577114 495436
rect 577332 495424 577366 495474
rect 577584 494292 577630 495436
rect 577698 495392 577744 495474
rect 562120 494221 567614 494277
rect 562120 494161 562222 494221
rect 562282 494161 562342 494221
rect 562402 494161 562462 494221
rect 562522 494161 562582 494221
rect 562642 494161 562702 494221
rect 562762 494161 562822 494221
rect 562882 494161 562942 494221
rect 563002 494161 563062 494221
rect 563122 494161 563182 494221
rect 563242 494161 563302 494221
rect 563362 494161 563422 494221
rect 563482 494161 563542 494221
rect 563602 494161 563662 494221
rect 563722 494161 563782 494221
rect 563842 494161 563902 494221
rect 563962 494161 564022 494221
rect 564082 494161 564142 494221
rect 564202 494161 564262 494221
rect 564322 494161 564382 494221
rect 564442 494161 564502 494221
rect 564562 494161 564622 494221
rect 564682 494161 564742 494221
rect 564802 494161 564862 494221
rect 564922 494161 564982 494221
rect 565042 494161 565102 494221
rect 565162 494161 565222 494221
rect 565282 494161 565342 494221
rect 565402 494161 565462 494221
rect 565522 494161 565582 494221
rect 565642 494161 565702 494221
rect 565762 494161 565822 494221
rect 565882 494161 565942 494221
rect 566002 494161 566062 494221
rect 566122 494161 566182 494221
rect 566242 494161 566302 494221
rect 566362 494161 566422 494221
rect 566482 494161 566542 494221
rect 566602 494161 566662 494221
rect 566722 494161 566782 494221
rect 566842 494161 566902 494221
rect 566962 494161 567022 494221
rect 567082 494161 567142 494221
rect 567202 494161 567262 494221
rect 567322 494161 567382 494221
rect 567442 494161 567502 494221
rect 567562 494161 567614 494221
rect 562120 494101 567614 494161
rect 562120 494041 562222 494101
rect 562282 494041 562342 494101
rect 562402 494041 562462 494101
rect 562522 494041 562582 494101
rect 562642 494041 562702 494101
rect 562762 494041 562822 494101
rect 562882 494041 562942 494101
rect 563002 494041 563062 494101
rect 563122 494041 563182 494101
rect 563242 494041 563302 494101
rect 563362 494041 563422 494101
rect 563482 494041 563542 494101
rect 563602 494041 563662 494101
rect 563722 494041 563782 494101
rect 563842 494041 563902 494101
rect 563962 494041 564022 494101
rect 564082 494041 564142 494101
rect 564202 494041 564262 494101
rect 564322 494041 564382 494101
rect 564442 494041 564502 494101
rect 564562 494041 564622 494101
rect 564682 494041 564742 494101
rect 564802 494041 564862 494101
rect 564922 494041 564982 494101
rect 565042 494041 565102 494101
rect 565162 494041 565222 494101
rect 565282 494041 565342 494101
rect 565402 494041 565462 494101
rect 565522 494041 565582 494101
rect 565642 494041 565702 494101
rect 565762 494041 565822 494101
rect 565882 494041 565942 494101
rect 566002 494041 566062 494101
rect 566122 494041 566182 494101
rect 566242 494041 566302 494101
rect 566362 494041 566422 494101
rect 566482 494041 566542 494101
rect 566602 494041 566662 494101
rect 566722 494041 566782 494101
rect 566842 494041 566902 494101
rect 566962 494041 567022 494101
rect 567082 494041 567142 494101
rect 567202 494041 567262 494101
rect 567322 494041 567382 494101
rect 567442 494041 567502 494101
rect 567562 494041 567614 494101
rect 562120 494002 567614 494041
rect 572280 494236 577774 494292
rect 572280 494176 572332 494236
rect 572392 494176 572452 494236
rect 572512 494176 572572 494236
rect 572632 494176 572692 494236
rect 572752 494176 572812 494236
rect 572872 494176 572932 494236
rect 572992 494176 573052 494236
rect 573112 494176 573172 494236
rect 573232 494176 573292 494236
rect 573352 494176 573412 494236
rect 573472 494176 573532 494236
rect 573592 494176 573652 494236
rect 573712 494176 573772 494236
rect 573832 494176 573892 494236
rect 573952 494176 574012 494236
rect 574072 494176 574132 494236
rect 574192 494176 574252 494236
rect 574312 494176 574372 494236
rect 574432 494176 574492 494236
rect 574552 494176 574612 494236
rect 574672 494176 574732 494236
rect 574792 494176 574852 494236
rect 574912 494176 574972 494236
rect 575032 494176 575092 494236
rect 575152 494176 575212 494236
rect 575272 494176 575332 494236
rect 575392 494176 575452 494236
rect 575512 494176 575572 494236
rect 575632 494176 575692 494236
rect 575752 494176 575812 494236
rect 575872 494176 575932 494236
rect 575992 494176 576052 494236
rect 576112 494176 576172 494236
rect 576232 494176 576292 494236
rect 576352 494176 576412 494236
rect 576472 494176 576532 494236
rect 576592 494176 576652 494236
rect 576712 494176 576772 494236
rect 576832 494176 576892 494236
rect 576952 494176 577012 494236
rect 577072 494176 577132 494236
rect 577192 494176 577252 494236
rect 577312 494176 577372 494236
rect 577432 494176 577492 494236
rect 577552 494176 577612 494236
rect 577672 494176 577774 494236
rect 572280 494116 577774 494176
rect 572280 494056 572332 494116
rect 572392 494056 572452 494116
rect 572512 494056 572572 494116
rect 572632 494056 572692 494116
rect 572752 494056 572812 494116
rect 572872 494056 572932 494116
rect 572992 494056 573052 494116
rect 573112 494056 573172 494116
rect 573232 494056 573292 494116
rect 573352 494056 573412 494116
rect 573472 494056 573532 494116
rect 573592 494056 573652 494116
rect 573712 494056 573772 494116
rect 573832 494056 573892 494116
rect 573952 494056 574012 494116
rect 574072 494056 574132 494116
rect 574192 494056 574252 494116
rect 574312 494056 574372 494116
rect 574432 494056 574492 494116
rect 574552 494056 574612 494116
rect 574672 494056 574732 494116
rect 574792 494056 574852 494116
rect 574912 494056 574972 494116
rect 575032 494056 575092 494116
rect 575152 494056 575212 494116
rect 575272 494056 575332 494116
rect 575392 494056 575452 494116
rect 575512 494056 575572 494116
rect 575632 494056 575692 494116
rect 575752 494056 575812 494116
rect 575872 494056 575932 494116
rect 575992 494056 576052 494116
rect 576112 494056 576172 494116
rect 576232 494056 576292 494116
rect 576352 494056 576412 494116
rect 576472 494056 576532 494116
rect 576592 494056 576652 494116
rect 576712 494056 576772 494116
rect 576832 494056 576892 494116
rect 576952 494056 577012 494116
rect 577072 494056 577132 494116
rect 577192 494056 577252 494116
rect 577312 494056 577372 494116
rect 577432 494056 577492 494116
rect 577552 494056 577612 494116
rect 577672 494056 577774 494116
rect 572280 494017 577774 494056
rect 562150 455440 567584 455473
rect 562150 455360 562480 455440
rect 562560 455360 562640 455440
rect 562720 455360 562800 455440
rect 562880 455360 562960 455440
rect 563040 455360 563120 455440
rect 563200 455360 563280 455440
rect 563360 455360 563440 455440
rect 563520 455360 563600 455440
rect 563680 455360 563760 455440
rect 563840 455360 563920 455440
rect 564000 455360 564080 455440
rect 564160 455360 564240 455440
rect 564320 455360 564400 455440
rect 564480 455360 564560 455440
rect 564640 455360 564720 455440
rect 564800 455360 564880 455440
rect 564960 455360 565040 455440
rect 565120 455360 565200 455440
rect 565280 455360 565360 455440
rect 565440 455360 565520 455440
rect 565600 455360 565680 455440
rect 565760 455360 565840 455440
rect 565920 455360 566000 455440
rect 566080 455360 566160 455440
rect 566240 455360 566320 455440
rect 566400 455360 566480 455440
rect 566560 455360 566640 455440
rect 566720 455360 566800 455440
rect 566880 455360 566960 455440
rect 567040 455360 567120 455440
rect 567200 455360 567280 455440
rect 567360 455360 567584 455440
rect 562150 455280 567584 455360
rect 562150 455200 562480 455280
rect 562560 455200 562640 455280
rect 562720 455200 562800 455280
rect 562880 455200 562960 455280
rect 563040 455200 563120 455280
rect 563200 455200 563280 455280
rect 563360 455200 563440 455280
rect 563520 455200 563600 455280
rect 563680 455200 563760 455280
rect 563840 455200 563920 455280
rect 564000 455200 564080 455280
rect 564160 455200 564240 455280
rect 564320 455200 564400 455280
rect 564480 455200 564560 455280
rect 564640 455200 564720 455280
rect 564800 455200 564880 455280
rect 564960 455200 565040 455280
rect 565120 455200 565200 455280
rect 565280 455200 565360 455280
rect 565440 455200 565520 455280
rect 565600 455200 565680 455280
rect 565760 455200 565840 455280
rect 565920 455200 566000 455280
rect 566080 455200 566160 455280
rect 566240 455200 566320 455280
rect 566400 455200 566480 455280
rect 566560 455200 566640 455280
rect 566720 455200 566800 455280
rect 566880 455200 566960 455280
rect 567040 455200 567120 455280
rect 567200 455200 567280 455280
rect 567360 455200 567584 455280
rect 562150 455172 567584 455200
rect 562150 454061 562196 455172
rect 562522 455100 562568 455172
rect 563038 455100 563084 455172
rect 563554 455100 563600 455172
rect 564070 455100 564116 455172
rect 564586 455100 564632 455172
rect 565102 455100 565148 455172
rect 565618 455100 565664 455172
rect 566134 455100 566180 455172
rect 566650 455100 566696 455172
rect 567166 455100 567212 455172
rect 562264 453975 562310 455100
rect 562780 453975 562826 455100
rect 563296 453975 563342 455100
rect 563812 453975 563858 455100
rect 564328 453975 564374 455100
rect 564844 453975 564890 455100
rect 565360 453975 565406 455100
rect 565876 453975 565922 455100
rect 566392 453975 566438 455100
rect 566908 453975 566954 455100
rect 567424 453975 567470 455100
rect 567538 454073 567584 455172
rect 572310 455440 577744 455473
rect 572310 455360 572640 455440
rect 572720 455360 572800 455440
rect 572880 455360 572960 455440
rect 573040 455360 573120 455440
rect 573200 455360 573280 455440
rect 573360 455360 573440 455440
rect 573520 455360 573600 455440
rect 573680 455360 573760 455440
rect 573840 455360 573920 455440
rect 574000 455360 574080 455440
rect 574160 455360 574240 455440
rect 574320 455360 574400 455440
rect 574480 455360 574560 455440
rect 574640 455360 574720 455440
rect 574800 455360 574880 455440
rect 574960 455360 575040 455440
rect 575120 455360 575200 455440
rect 575280 455360 575360 455440
rect 575440 455360 575520 455440
rect 575600 455360 575680 455440
rect 575760 455360 575840 455440
rect 575920 455360 576000 455440
rect 576080 455360 576160 455440
rect 576240 455360 576320 455440
rect 576400 455360 576480 455440
rect 576560 455360 576640 455440
rect 576720 455360 576800 455440
rect 576880 455360 576960 455440
rect 577040 455360 577120 455440
rect 577200 455360 577280 455440
rect 577360 455360 577440 455440
rect 577520 455360 577744 455440
rect 572310 455280 577744 455360
rect 572310 455200 572640 455280
rect 572720 455200 572800 455280
rect 572880 455200 572960 455280
rect 573040 455200 573120 455280
rect 573200 455200 573280 455280
rect 573360 455200 573440 455280
rect 573520 455200 573600 455280
rect 573680 455200 573760 455280
rect 573840 455200 573920 455280
rect 574000 455200 574080 455280
rect 574160 455200 574240 455280
rect 574320 455200 574400 455280
rect 574480 455200 574560 455280
rect 574640 455200 574720 455280
rect 574800 455200 574880 455280
rect 574960 455200 575040 455280
rect 575120 455200 575200 455280
rect 575280 455200 575360 455280
rect 575440 455200 575520 455280
rect 575600 455200 575680 455280
rect 575760 455200 575840 455280
rect 575920 455200 576000 455280
rect 576080 455200 576160 455280
rect 576240 455200 576320 455280
rect 576400 455200 576480 455280
rect 576560 455200 576640 455280
rect 576720 455200 576800 455280
rect 576880 455200 576960 455280
rect 577040 455200 577120 455280
rect 577200 455200 577280 455280
rect 577360 455200 577440 455280
rect 577520 455200 577744 455280
rect 572310 455172 577744 455200
rect 572310 455090 572356 455172
rect 572424 453990 572470 455134
rect 572688 455122 572722 455172
rect 572940 453990 572986 455134
rect 573204 455122 573238 455172
rect 573456 453990 573502 455134
rect 573720 455122 573754 455172
rect 573972 453990 574018 455134
rect 574236 455122 574270 455172
rect 574488 453990 574534 455134
rect 574752 455122 574786 455172
rect 575004 453990 575050 455134
rect 575268 455122 575302 455172
rect 575520 453990 575566 455134
rect 575784 455122 575818 455172
rect 576036 453990 576082 455134
rect 576300 455122 576334 455172
rect 576552 453990 576598 455134
rect 576816 455122 576850 455172
rect 577068 453990 577114 455134
rect 577332 455122 577366 455172
rect 577584 453990 577630 455134
rect 577698 455090 577744 455172
rect 562120 453919 567614 453975
rect 562120 453859 562222 453919
rect 562282 453859 562342 453919
rect 562402 453859 562462 453919
rect 562522 453859 562582 453919
rect 562642 453859 562702 453919
rect 562762 453859 562822 453919
rect 562882 453859 562942 453919
rect 563002 453859 563062 453919
rect 563122 453859 563182 453919
rect 563242 453859 563302 453919
rect 563362 453859 563422 453919
rect 563482 453859 563542 453919
rect 563602 453859 563662 453919
rect 563722 453859 563782 453919
rect 563842 453859 563902 453919
rect 563962 453859 564022 453919
rect 564082 453859 564142 453919
rect 564202 453859 564262 453919
rect 564322 453859 564382 453919
rect 564442 453859 564502 453919
rect 564562 453859 564622 453919
rect 564682 453859 564742 453919
rect 564802 453859 564862 453919
rect 564922 453859 564982 453919
rect 565042 453859 565102 453919
rect 565162 453859 565222 453919
rect 565282 453859 565342 453919
rect 565402 453859 565462 453919
rect 565522 453859 565582 453919
rect 565642 453859 565702 453919
rect 565762 453859 565822 453919
rect 565882 453859 565942 453919
rect 566002 453859 566062 453919
rect 566122 453859 566182 453919
rect 566242 453859 566302 453919
rect 566362 453859 566422 453919
rect 566482 453859 566542 453919
rect 566602 453859 566662 453919
rect 566722 453859 566782 453919
rect 566842 453859 566902 453919
rect 566962 453859 567022 453919
rect 567082 453859 567142 453919
rect 567202 453859 567262 453919
rect 567322 453859 567382 453919
rect 567442 453859 567502 453919
rect 567562 453859 567614 453919
rect 562120 453799 567614 453859
rect 562120 453739 562222 453799
rect 562282 453739 562342 453799
rect 562402 453739 562462 453799
rect 562522 453739 562582 453799
rect 562642 453739 562702 453799
rect 562762 453739 562822 453799
rect 562882 453739 562942 453799
rect 563002 453739 563062 453799
rect 563122 453739 563182 453799
rect 563242 453739 563302 453799
rect 563362 453739 563422 453799
rect 563482 453739 563542 453799
rect 563602 453739 563662 453799
rect 563722 453739 563782 453799
rect 563842 453739 563902 453799
rect 563962 453739 564022 453799
rect 564082 453739 564142 453799
rect 564202 453739 564262 453799
rect 564322 453739 564382 453799
rect 564442 453739 564502 453799
rect 564562 453739 564622 453799
rect 564682 453739 564742 453799
rect 564802 453739 564862 453799
rect 564922 453739 564982 453799
rect 565042 453739 565102 453799
rect 565162 453739 565222 453799
rect 565282 453739 565342 453799
rect 565402 453739 565462 453799
rect 565522 453739 565582 453799
rect 565642 453739 565702 453799
rect 565762 453739 565822 453799
rect 565882 453739 565942 453799
rect 566002 453739 566062 453799
rect 566122 453739 566182 453799
rect 566242 453739 566302 453799
rect 566362 453739 566422 453799
rect 566482 453739 566542 453799
rect 566602 453739 566662 453799
rect 566722 453739 566782 453799
rect 566842 453739 566902 453799
rect 566962 453739 567022 453799
rect 567082 453739 567142 453799
rect 567202 453739 567262 453799
rect 567322 453739 567382 453799
rect 567442 453739 567502 453799
rect 567562 453739 567614 453799
rect 562120 453700 567614 453739
rect 572280 453934 577774 453990
rect 572280 453874 572332 453934
rect 572392 453874 572452 453934
rect 572512 453874 572572 453934
rect 572632 453874 572692 453934
rect 572752 453874 572812 453934
rect 572872 453874 572932 453934
rect 572992 453874 573052 453934
rect 573112 453874 573172 453934
rect 573232 453874 573292 453934
rect 573352 453874 573412 453934
rect 573472 453874 573532 453934
rect 573592 453874 573652 453934
rect 573712 453874 573772 453934
rect 573832 453874 573892 453934
rect 573952 453874 574012 453934
rect 574072 453874 574132 453934
rect 574192 453874 574252 453934
rect 574312 453874 574372 453934
rect 574432 453874 574492 453934
rect 574552 453874 574612 453934
rect 574672 453874 574732 453934
rect 574792 453874 574852 453934
rect 574912 453874 574972 453934
rect 575032 453874 575092 453934
rect 575152 453874 575212 453934
rect 575272 453874 575332 453934
rect 575392 453874 575452 453934
rect 575512 453874 575572 453934
rect 575632 453874 575692 453934
rect 575752 453874 575812 453934
rect 575872 453874 575932 453934
rect 575992 453874 576052 453934
rect 576112 453874 576172 453934
rect 576232 453874 576292 453934
rect 576352 453874 576412 453934
rect 576472 453874 576532 453934
rect 576592 453874 576652 453934
rect 576712 453874 576772 453934
rect 576832 453874 576892 453934
rect 576952 453874 577012 453934
rect 577072 453874 577132 453934
rect 577192 453874 577252 453934
rect 577312 453874 577372 453934
rect 577432 453874 577492 453934
rect 577552 453874 577612 453934
rect 577672 453874 577774 453934
rect 572280 453814 577774 453874
rect 572280 453754 572332 453814
rect 572392 453754 572452 453814
rect 572512 453754 572572 453814
rect 572632 453754 572692 453814
rect 572752 453754 572812 453814
rect 572872 453754 572932 453814
rect 572992 453754 573052 453814
rect 573112 453754 573172 453814
rect 573232 453754 573292 453814
rect 573352 453754 573412 453814
rect 573472 453754 573532 453814
rect 573592 453754 573652 453814
rect 573712 453754 573772 453814
rect 573832 453754 573892 453814
rect 573952 453754 574012 453814
rect 574072 453754 574132 453814
rect 574192 453754 574252 453814
rect 574312 453754 574372 453814
rect 574432 453754 574492 453814
rect 574552 453754 574612 453814
rect 574672 453754 574732 453814
rect 574792 453754 574852 453814
rect 574912 453754 574972 453814
rect 575032 453754 575092 453814
rect 575152 453754 575212 453814
rect 575272 453754 575332 453814
rect 575392 453754 575452 453814
rect 575512 453754 575572 453814
rect 575632 453754 575692 453814
rect 575752 453754 575812 453814
rect 575872 453754 575932 453814
rect 575992 453754 576052 453814
rect 576112 453754 576172 453814
rect 576232 453754 576292 453814
rect 576352 453754 576412 453814
rect 576472 453754 576532 453814
rect 576592 453754 576652 453814
rect 576712 453754 576772 453814
rect 576832 453754 576892 453814
rect 576952 453754 577012 453814
rect 577072 453754 577132 453814
rect 577192 453754 577252 453814
rect 577312 453754 577372 453814
rect 577432 453754 577492 453814
rect 577552 453754 577612 453814
rect 577672 453754 577774 453814
rect 572280 453715 577774 453754
<< via1 >>
rect 562480 495662 562560 495742
rect 562640 495662 562720 495742
rect 562800 495662 562880 495742
rect 562960 495662 563040 495742
rect 563120 495662 563200 495742
rect 563280 495662 563360 495742
rect 563440 495662 563520 495742
rect 563600 495662 563680 495742
rect 563760 495662 563840 495742
rect 563920 495662 564000 495742
rect 564080 495662 564160 495742
rect 564240 495662 564320 495742
rect 564400 495662 564480 495742
rect 564560 495662 564640 495742
rect 564720 495662 564800 495742
rect 564880 495662 564960 495742
rect 565040 495662 565120 495742
rect 565200 495662 565280 495742
rect 565360 495662 565440 495742
rect 565520 495662 565600 495742
rect 565680 495662 565760 495742
rect 565840 495662 565920 495742
rect 566000 495662 566080 495742
rect 566160 495662 566240 495742
rect 566320 495662 566400 495742
rect 566480 495662 566560 495742
rect 566640 495662 566720 495742
rect 566800 495662 566880 495742
rect 566960 495662 567040 495742
rect 567120 495662 567200 495742
rect 567280 495662 567360 495742
rect 562480 495502 562560 495582
rect 562640 495502 562720 495582
rect 562800 495502 562880 495582
rect 562960 495502 563040 495582
rect 563120 495502 563200 495582
rect 563280 495502 563360 495582
rect 563440 495502 563520 495582
rect 563600 495502 563680 495582
rect 563760 495502 563840 495582
rect 563920 495502 564000 495582
rect 564080 495502 564160 495582
rect 564240 495502 564320 495582
rect 564400 495502 564480 495582
rect 564560 495502 564640 495582
rect 564720 495502 564800 495582
rect 564880 495502 564960 495582
rect 565040 495502 565120 495582
rect 565200 495502 565280 495582
rect 565360 495502 565440 495582
rect 565520 495502 565600 495582
rect 565680 495502 565760 495582
rect 565840 495502 565920 495582
rect 566000 495502 566080 495582
rect 566160 495502 566240 495582
rect 566320 495502 566400 495582
rect 566480 495502 566560 495582
rect 566640 495502 566720 495582
rect 566800 495502 566880 495582
rect 566960 495502 567040 495582
rect 567120 495502 567200 495582
rect 567280 495502 567360 495582
rect 572640 495662 572720 495742
rect 572800 495662 572880 495742
rect 572960 495662 573040 495742
rect 573120 495662 573200 495742
rect 573280 495662 573360 495742
rect 573440 495662 573520 495742
rect 573600 495662 573680 495742
rect 573760 495662 573840 495742
rect 573920 495662 574000 495742
rect 574080 495662 574160 495742
rect 574240 495662 574320 495742
rect 574400 495662 574480 495742
rect 574560 495662 574640 495742
rect 574720 495662 574800 495742
rect 574880 495662 574960 495742
rect 575040 495662 575120 495742
rect 575200 495662 575280 495742
rect 575360 495662 575440 495742
rect 575520 495662 575600 495742
rect 575680 495662 575760 495742
rect 575840 495662 575920 495742
rect 576000 495662 576080 495742
rect 576160 495662 576240 495742
rect 576320 495662 576400 495742
rect 576480 495662 576560 495742
rect 576640 495662 576720 495742
rect 576800 495662 576880 495742
rect 576960 495662 577040 495742
rect 577120 495662 577200 495742
rect 577280 495662 577360 495742
rect 577440 495662 577520 495742
rect 572640 495502 572720 495582
rect 572800 495502 572880 495582
rect 572960 495502 573040 495582
rect 573120 495502 573200 495582
rect 573280 495502 573360 495582
rect 573440 495502 573520 495582
rect 573600 495502 573680 495582
rect 573760 495502 573840 495582
rect 573920 495502 574000 495582
rect 574080 495502 574160 495582
rect 574240 495502 574320 495582
rect 574400 495502 574480 495582
rect 574560 495502 574640 495582
rect 574720 495502 574800 495582
rect 574880 495502 574960 495582
rect 575040 495502 575120 495582
rect 575200 495502 575280 495582
rect 575360 495502 575440 495582
rect 575520 495502 575600 495582
rect 575680 495502 575760 495582
rect 575840 495502 575920 495582
rect 576000 495502 576080 495582
rect 576160 495502 576240 495582
rect 576320 495502 576400 495582
rect 576480 495502 576560 495582
rect 576640 495502 576720 495582
rect 576800 495502 576880 495582
rect 576960 495502 577040 495582
rect 577120 495502 577200 495582
rect 577280 495502 577360 495582
rect 577440 495502 577520 495582
rect 562222 494161 562282 494221
rect 562342 494161 562402 494221
rect 562462 494161 562522 494221
rect 562582 494161 562642 494221
rect 562702 494161 562762 494221
rect 562822 494161 562882 494221
rect 562942 494161 563002 494221
rect 563062 494161 563122 494221
rect 563182 494161 563242 494221
rect 563302 494161 563362 494221
rect 563422 494161 563482 494221
rect 563542 494161 563602 494221
rect 563662 494161 563722 494221
rect 563782 494161 563842 494221
rect 563902 494161 563962 494221
rect 564022 494161 564082 494221
rect 564142 494161 564202 494221
rect 564262 494161 564322 494221
rect 564382 494161 564442 494221
rect 564502 494161 564562 494221
rect 564622 494161 564682 494221
rect 564742 494161 564802 494221
rect 564862 494161 564922 494221
rect 564982 494161 565042 494221
rect 565102 494161 565162 494221
rect 565222 494161 565282 494221
rect 565342 494161 565402 494221
rect 565462 494161 565522 494221
rect 565582 494161 565642 494221
rect 565702 494161 565762 494221
rect 565822 494161 565882 494221
rect 565942 494161 566002 494221
rect 566062 494161 566122 494221
rect 566182 494161 566242 494221
rect 566302 494161 566362 494221
rect 566422 494161 566482 494221
rect 566542 494161 566602 494221
rect 566662 494161 566722 494221
rect 566782 494161 566842 494221
rect 566902 494161 566962 494221
rect 567022 494161 567082 494221
rect 567142 494161 567202 494221
rect 567262 494161 567322 494221
rect 567382 494161 567442 494221
rect 567502 494161 567562 494221
rect 562222 494041 562282 494101
rect 562342 494041 562402 494101
rect 562462 494041 562522 494101
rect 562582 494041 562642 494101
rect 562702 494041 562762 494101
rect 562822 494041 562882 494101
rect 562942 494041 563002 494101
rect 563062 494041 563122 494101
rect 563182 494041 563242 494101
rect 563302 494041 563362 494101
rect 563422 494041 563482 494101
rect 563542 494041 563602 494101
rect 563662 494041 563722 494101
rect 563782 494041 563842 494101
rect 563902 494041 563962 494101
rect 564022 494041 564082 494101
rect 564142 494041 564202 494101
rect 564262 494041 564322 494101
rect 564382 494041 564442 494101
rect 564502 494041 564562 494101
rect 564622 494041 564682 494101
rect 564742 494041 564802 494101
rect 564862 494041 564922 494101
rect 564982 494041 565042 494101
rect 565102 494041 565162 494101
rect 565222 494041 565282 494101
rect 565342 494041 565402 494101
rect 565462 494041 565522 494101
rect 565582 494041 565642 494101
rect 565702 494041 565762 494101
rect 565822 494041 565882 494101
rect 565942 494041 566002 494101
rect 566062 494041 566122 494101
rect 566182 494041 566242 494101
rect 566302 494041 566362 494101
rect 566422 494041 566482 494101
rect 566542 494041 566602 494101
rect 566662 494041 566722 494101
rect 566782 494041 566842 494101
rect 566902 494041 566962 494101
rect 567022 494041 567082 494101
rect 567142 494041 567202 494101
rect 567262 494041 567322 494101
rect 567382 494041 567442 494101
rect 567502 494041 567562 494101
rect 572332 494176 572392 494236
rect 572452 494176 572512 494236
rect 572572 494176 572632 494236
rect 572692 494176 572752 494236
rect 572812 494176 572872 494236
rect 572932 494176 572992 494236
rect 573052 494176 573112 494236
rect 573172 494176 573232 494236
rect 573292 494176 573352 494236
rect 573412 494176 573472 494236
rect 573532 494176 573592 494236
rect 573652 494176 573712 494236
rect 573772 494176 573832 494236
rect 573892 494176 573952 494236
rect 574012 494176 574072 494236
rect 574132 494176 574192 494236
rect 574252 494176 574312 494236
rect 574372 494176 574432 494236
rect 574492 494176 574552 494236
rect 574612 494176 574672 494236
rect 574732 494176 574792 494236
rect 574852 494176 574912 494236
rect 574972 494176 575032 494236
rect 575092 494176 575152 494236
rect 575212 494176 575272 494236
rect 575332 494176 575392 494236
rect 575452 494176 575512 494236
rect 575572 494176 575632 494236
rect 575692 494176 575752 494236
rect 575812 494176 575872 494236
rect 575932 494176 575992 494236
rect 576052 494176 576112 494236
rect 576172 494176 576232 494236
rect 576292 494176 576352 494236
rect 576412 494176 576472 494236
rect 576532 494176 576592 494236
rect 576652 494176 576712 494236
rect 576772 494176 576832 494236
rect 576892 494176 576952 494236
rect 577012 494176 577072 494236
rect 577132 494176 577192 494236
rect 577252 494176 577312 494236
rect 577372 494176 577432 494236
rect 577492 494176 577552 494236
rect 577612 494176 577672 494236
rect 572332 494056 572392 494116
rect 572452 494056 572512 494116
rect 572572 494056 572632 494116
rect 572692 494056 572752 494116
rect 572812 494056 572872 494116
rect 572932 494056 572992 494116
rect 573052 494056 573112 494116
rect 573172 494056 573232 494116
rect 573292 494056 573352 494116
rect 573412 494056 573472 494116
rect 573532 494056 573592 494116
rect 573652 494056 573712 494116
rect 573772 494056 573832 494116
rect 573892 494056 573952 494116
rect 574012 494056 574072 494116
rect 574132 494056 574192 494116
rect 574252 494056 574312 494116
rect 574372 494056 574432 494116
rect 574492 494056 574552 494116
rect 574612 494056 574672 494116
rect 574732 494056 574792 494116
rect 574852 494056 574912 494116
rect 574972 494056 575032 494116
rect 575092 494056 575152 494116
rect 575212 494056 575272 494116
rect 575332 494056 575392 494116
rect 575452 494056 575512 494116
rect 575572 494056 575632 494116
rect 575692 494056 575752 494116
rect 575812 494056 575872 494116
rect 575932 494056 575992 494116
rect 576052 494056 576112 494116
rect 576172 494056 576232 494116
rect 576292 494056 576352 494116
rect 576412 494056 576472 494116
rect 576532 494056 576592 494116
rect 576652 494056 576712 494116
rect 576772 494056 576832 494116
rect 576892 494056 576952 494116
rect 577012 494056 577072 494116
rect 577132 494056 577192 494116
rect 577252 494056 577312 494116
rect 577372 494056 577432 494116
rect 577492 494056 577552 494116
rect 577612 494056 577672 494116
rect 562480 455360 562560 455440
rect 562640 455360 562720 455440
rect 562800 455360 562880 455440
rect 562960 455360 563040 455440
rect 563120 455360 563200 455440
rect 563280 455360 563360 455440
rect 563440 455360 563520 455440
rect 563600 455360 563680 455440
rect 563760 455360 563840 455440
rect 563920 455360 564000 455440
rect 564080 455360 564160 455440
rect 564240 455360 564320 455440
rect 564400 455360 564480 455440
rect 564560 455360 564640 455440
rect 564720 455360 564800 455440
rect 564880 455360 564960 455440
rect 565040 455360 565120 455440
rect 565200 455360 565280 455440
rect 565360 455360 565440 455440
rect 565520 455360 565600 455440
rect 565680 455360 565760 455440
rect 565840 455360 565920 455440
rect 566000 455360 566080 455440
rect 566160 455360 566240 455440
rect 566320 455360 566400 455440
rect 566480 455360 566560 455440
rect 566640 455360 566720 455440
rect 566800 455360 566880 455440
rect 566960 455360 567040 455440
rect 567120 455360 567200 455440
rect 567280 455360 567360 455440
rect 562480 455200 562560 455280
rect 562640 455200 562720 455280
rect 562800 455200 562880 455280
rect 562960 455200 563040 455280
rect 563120 455200 563200 455280
rect 563280 455200 563360 455280
rect 563440 455200 563520 455280
rect 563600 455200 563680 455280
rect 563760 455200 563840 455280
rect 563920 455200 564000 455280
rect 564080 455200 564160 455280
rect 564240 455200 564320 455280
rect 564400 455200 564480 455280
rect 564560 455200 564640 455280
rect 564720 455200 564800 455280
rect 564880 455200 564960 455280
rect 565040 455200 565120 455280
rect 565200 455200 565280 455280
rect 565360 455200 565440 455280
rect 565520 455200 565600 455280
rect 565680 455200 565760 455280
rect 565840 455200 565920 455280
rect 566000 455200 566080 455280
rect 566160 455200 566240 455280
rect 566320 455200 566400 455280
rect 566480 455200 566560 455280
rect 566640 455200 566720 455280
rect 566800 455200 566880 455280
rect 566960 455200 567040 455280
rect 567120 455200 567200 455280
rect 567280 455200 567360 455280
rect 572640 455360 572720 455440
rect 572800 455360 572880 455440
rect 572960 455360 573040 455440
rect 573120 455360 573200 455440
rect 573280 455360 573360 455440
rect 573440 455360 573520 455440
rect 573600 455360 573680 455440
rect 573760 455360 573840 455440
rect 573920 455360 574000 455440
rect 574080 455360 574160 455440
rect 574240 455360 574320 455440
rect 574400 455360 574480 455440
rect 574560 455360 574640 455440
rect 574720 455360 574800 455440
rect 574880 455360 574960 455440
rect 575040 455360 575120 455440
rect 575200 455360 575280 455440
rect 575360 455360 575440 455440
rect 575520 455360 575600 455440
rect 575680 455360 575760 455440
rect 575840 455360 575920 455440
rect 576000 455360 576080 455440
rect 576160 455360 576240 455440
rect 576320 455360 576400 455440
rect 576480 455360 576560 455440
rect 576640 455360 576720 455440
rect 576800 455360 576880 455440
rect 576960 455360 577040 455440
rect 577120 455360 577200 455440
rect 577280 455360 577360 455440
rect 577440 455360 577520 455440
rect 572640 455200 572720 455280
rect 572800 455200 572880 455280
rect 572960 455200 573040 455280
rect 573120 455200 573200 455280
rect 573280 455200 573360 455280
rect 573440 455200 573520 455280
rect 573600 455200 573680 455280
rect 573760 455200 573840 455280
rect 573920 455200 574000 455280
rect 574080 455200 574160 455280
rect 574240 455200 574320 455280
rect 574400 455200 574480 455280
rect 574560 455200 574640 455280
rect 574720 455200 574800 455280
rect 574880 455200 574960 455280
rect 575040 455200 575120 455280
rect 575200 455200 575280 455280
rect 575360 455200 575440 455280
rect 575520 455200 575600 455280
rect 575680 455200 575760 455280
rect 575840 455200 575920 455280
rect 576000 455200 576080 455280
rect 576160 455200 576240 455280
rect 576320 455200 576400 455280
rect 576480 455200 576560 455280
rect 576640 455200 576720 455280
rect 576800 455200 576880 455280
rect 576960 455200 577040 455280
rect 577120 455200 577200 455280
rect 577280 455200 577360 455280
rect 577440 455200 577520 455280
rect 562222 453859 562282 453919
rect 562342 453859 562402 453919
rect 562462 453859 562522 453919
rect 562582 453859 562642 453919
rect 562702 453859 562762 453919
rect 562822 453859 562882 453919
rect 562942 453859 563002 453919
rect 563062 453859 563122 453919
rect 563182 453859 563242 453919
rect 563302 453859 563362 453919
rect 563422 453859 563482 453919
rect 563542 453859 563602 453919
rect 563662 453859 563722 453919
rect 563782 453859 563842 453919
rect 563902 453859 563962 453919
rect 564022 453859 564082 453919
rect 564142 453859 564202 453919
rect 564262 453859 564322 453919
rect 564382 453859 564442 453919
rect 564502 453859 564562 453919
rect 564622 453859 564682 453919
rect 564742 453859 564802 453919
rect 564862 453859 564922 453919
rect 564982 453859 565042 453919
rect 565102 453859 565162 453919
rect 565222 453859 565282 453919
rect 565342 453859 565402 453919
rect 565462 453859 565522 453919
rect 565582 453859 565642 453919
rect 565702 453859 565762 453919
rect 565822 453859 565882 453919
rect 565942 453859 566002 453919
rect 566062 453859 566122 453919
rect 566182 453859 566242 453919
rect 566302 453859 566362 453919
rect 566422 453859 566482 453919
rect 566542 453859 566602 453919
rect 566662 453859 566722 453919
rect 566782 453859 566842 453919
rect 566902 453859 566962 453919
rect 567022 453859 567082 453919
rect 567142 453859 567202 453919
rect 567262 453859 567322 453919
rect 567382 453859 567442 453919
rect 567502 453859 567562 453919
rect 562222 453739 562282 453799
rect 562342 453739 562402 453799
rect 562462 453739 562522 453799
rect 562582 453739 562642 453799
rect 562702 453739 562762 453799
rect 562822 453739 562882 453799
rect 562942 453739 563002 453799
rect 563062 453739 563122 453799
rect 563182 453739 563242 453799
rect 563302 453739 563362 453799
rect 563422 453739 563482 453799
rect 563542 453739 563602 453799
rect 563662 453739 563722 453799
rect 563782 453739 563842 453799
rect 563902 453739 563962 453799
rect 564022 453739 564082 453799
rect 564142 453739 564202 453799
rect 564262 453739 564322 453799
rect 564382 453739 564442 453799
rect 564502 453739 564562 453799
rect 564622 453739 564682 453799
rect 564742 453739 564802 453799
rect 564862 453739 564922 453799
rect 564982 453739 565042 453799
rect 565102 453739 565162 453799
rect 565222 453739 565282 453799
rect 565342 453739 565402 453799
rect 565462 453739 565522 453799
rect 565582 453739 565642 453799
rect 565702 453739 565762 453799
rect 565822 453739 565882 453799
rect 565942 453739 566002 453799
rect 566062 453739 566122 453799
rect 566182 453739 566242 453799
rect 566302 453739 566362 453799
rect 566422 453739 566482 453799
rect 566542 453739 566602 453799
rect 566662 453739 566722 453799
rect 566782 453739 566842 453799
rect 566902 453739 566962 453799
rect 567022 453739 567082 453799
rect 567142 453739 567202 453799
rect 567262 453739 567322 453799
rect 567382 453739 567442 453799
rect 567502 453739 567562 453799
rect 572332 453874 572392 453934
rect 572452 453874 572512 453934
rect 572572 453874 572632 453934
rect 572692 453874 572752 453934
rect 572812 453874 572872 453934
rect 572932 453874 572992 453934
rect 573052 453874 573112 453934
rect 573172 453874 573232 453934
rect 573292 453874 573352 453934
rect 573412 453874 573472 453934
rect 573532 453874 573592 453934
rect 573652 453874 573712 453934
rect 573772 453874 573832 453934
rect 573892 453874 573952 453934
rect 574012 453874 574072 453934
rect 574132 453874 574192 453934
rect 574252 453874 574312 453934
rect 574372 453874 574432 453934
rect 574492 453874 574552 453934
rect 574612 453874 574672 453934
rect 574732 453874 574792 453934
rect 574852 453874 574912 453934
rect 574972 453874 575032 453934
rect 575092 453874 575152 453934
rect 575212 453874 575272 453934
rect 575332 453874 575392 453934
rect 575452 453874 575512 453934
rect 575572 453874 575632 453934
rect 575692 453874 575752 453934
rect 575812 453874 575872 453934
rect 575932 453874 575992 453934
rect 576052 453874 576112 453934
rect 576172 453874 576232 453934
rect 576292 453874 576352 453934
rect 576412 453874 576472 453934
rect 576532 453874 576592 453934
rect 576652 453874 576712 453934
rect 576772 453874 576832 453934
rect 576892 453874 576952 453934
rect 577012 453874 577072 453934
rect 577132 453874 577192 453934
rect 577252 453874 577312 453934
rect 577372 453874 577432 453934
rect 577492 453874 577552 453934
rect 577612 453874 577672 453934
rect 572332 453754 572392 453814
rect 572452 453754 572512 453814
rect 572572 453754 572632 453814
rect 572692 453754 572752 453814
rect 572812 453754 572872 453814
rect 572932 453754 572992 453814
rect 573052 453754 573112 453814
rect 573172 453754 573232 453814
rect 573292 453754 573352 453814
rect 573412 453754 573472 453814
rect 573532 453754 573592 453814
rect 573652 453754 573712 453814
rect 573772 453754 573832 453814
rect 573892 453754 573952 453814
rect 574012 453754 574072 453814
rect 574132 453754 574192 453814
rect 574252 453754 574312 453814
rect 574372 453754 574432 453814
rect 574492 453754 574552 453814
rect 574612 453754 574672 453814
rect 574732 453754 574792 453814
rect 574852 453754 574912 453814
rect 574972 453754 575032 453814
rect 575092 453754 575152 453814
rect 575212 453754 575272 453814
rect 575332 453754 575392 453814
rect 575452 453754 575512 453814
rect 575572 453754 575632 453814
rect 575692 453754 575752 453814
rect 575812 453754 575872 453814
rect 575932 453754 575992 453814
rect 576052 453754 576112 453814
rect 576172 453754 576232 453814
rect 576292 453754 576352 453814
rect 576412 453754 576472 453814
rect 576532 453754 576592 453814
rect 576652 453754 576712 453814
rect 576772 453754 576832 453814
rect 576892 453754 576952 453814
rect 577012 453754 577072 453814
rect 577132 453754 577192 453814
rect 577252 453754 577312 453814
rect 577372 453754 577432 453814
rect 577492 453754 577552 453814
rect 577612 453754 577672 453814
<< metal2 >>
rect 562380 495742 567480 495822
rect 562380 495662 562480 495742
rect 562560 495662 562640 495742
rect 562720 495662 562800 495742
rect 562880 495662 562960 495742
rect 563040 495662 563120 495742
rect 563200 495662 563280 495742
rect 563360 495662 563440 495742
rect 563520 495662 563600 495742
rect 563680 495662 563760 495742
rect 563840 495662 563920 495742
rect 564000 495662 564080 495742
rect 564160 495662 564240 495742
rect 564320 495662 564400 495742
rect 564480 495662 564560 495742
rect 564640 495662 564720 495742
rect 564800 495662 564880 495742
rect 564960 495662 565040 495742
rect 565120 495662 565200 495742
rect 565280 495662 565360 495742
rect 565440 495662 565520 495742
rect 565600 495662 565680 495742
rect 565760 495662 565840 495742
rect 565920 495662 566000 495742
rect 566080 495662 566160 495742
rect 566240 495662 566320 495742
rect 566400 495662 566480 495742
rect 566560 495662 566640 495742
rect 566720 495662 566800 495742
rect 566880 495662 566960 495742
rect 567040 495662 567120 495742
rect 567200 495662 567280 495742
rect 567360 495662 567480 495742
rect 562380 495582 567480 495662
rect 562380 495502 562480 495582
rect 562560 495502 562640 495582
rect 562720 495502 562800 495582
rect 562880 495502 562960 495582
rect 563040 495502 563120 495582
rect 563200 495502 563280 495582
rect 563360 495502 563440 495582
rect 563520 495502 563600 495582
rect 563680 495502 563760 495582
rect 563840 495502 563920 495582
rect 564000 495502 564080 495582
rect 564160 495502 564240 495582
rect 564320 495502 564400 495582
rect 564480 495502 564560 495582
rect 564640 495502 564720 495582
rect 564800 495502 564880 495582
rect 564960 495502 565040 495582
rect 565120 495502 565200 495582
rect 565280 495502 565360 495582
rect 565440 495502 565520 495582
rect 565600 495502 565680 495582
rect 565760 495502 565840 495582
rect 565920 495502 566000 495582
rect 566080 495502 566160 495582
rect 566240 495502 566320 495582
rect 566400 495502 566480 495582
rect 566560 495502 566640 495582
rect 566720 495502 566800 495582
rect 566880 495502 566960 495582
rect 567040 495502 567120 495582
rect 567200 495502 567280 495582
rect 567360 495502 567480 495582
rect 562380 495462 567480 495502
rect 572540 495742 577640 495822
rect 572540 495662 572640 495742
rect 572720 495662 572800 495742
rect 572880 495662 572960 495742
rect 573040 495662 573120 495742
rect 573200 495662 573280 495742
rect 573360 495662 573440 495742
rect 573520 495662 573600 495742
rect 573680 495662 573760 495742
rect 573840 495662 573920 495742
rect 574000 495662 574080 495742
rect 574160 495662 574240 495742
rect 574320 495662 574400 495742
rect 574480 495662 574560 495742
rect 574640 495662 574720 495742
rect 574800 495662 574880 495742
rect 574960 495662 575040 495742
rect 575120 495662 575200 495742
rect 575280 495662 575360 495742
rect 575440 495662 575520 495742
rect 575600 495662 575680 495742
rect 575760 495662 575840 495742
rect 575920 495662 576000 495742
rect 576080 495662 576160 495742
rect 576240 495662 576320 495742
rect 576400 495662 576480 495742
rect 576560 495662 576640 495742
rect 576720 495662 576800 495742
rect 576880 495662 576960 495742
rect 577040 495662 577120 495742
rect 577200 495662 577280 495742
rect 577360 495662 577440 495742
rect 577520 495662 577640 495742
rect 572540 495582 577640 495662
rect 572540 495502 572640 495582
rect 572720 495502 572800 495582
rect 572880 495502 572960 495582
rect 573040 495502 573120 495582
rect 573200 495502 573280 495582
rect 573360 495502 573440 495582
rect 573520 495502 573600 495582
rect 573680 495502 573760 495582
rect 573840 495502 573920 495582
rect 574000 495502 574080 495582
rect 574160 495502 574240 495582
rect 574320 495502 574400 495582
rect 574480 495502 574560 495582
rect 574640 495502 574720 495582
rect 574800 495502 574880 495582
rect 574960 495502 575040 495582
rect 575120 495502 575200 495582
rect 575280 495502 575360 495582
rect 575440 495502 575520 495582
rect 575600 495502 575680 495582
rect 575760 495502 575840 495582
rect 575920 495502 576000 495582
rect 576080 495502 576160 495582
rect 576240 495502 576320 495582
rect 576400 495502 576480 495582
rect 576560 495502 576640 495582
rect 576720 495502 576800 495582
rect 576880 495502 576960 495582
rect 577040 495502 577120 495582
rect 577200 495502 577280 495582
rect 577360 495502 577440 495582
rect 577520 495502 577640 495582
rect 572540 495462 577640 495502
rect 562102 494221 567622 494281
rect 562102 494161 562222 494221
rect 562282 494161 562342 494221
rect 562402 494161 562462 494221
rect 562522 494161 562582 494221
rect 562642 494161 562702 494221
rect 562762 494161 562822 494221
rect 562882 494161 562942 494221
rect 563002 494161 563062 494221
rect 563122 494161 563182 494221
rect 563242 494161 563302 494221
rect 563362 494161 563422 494221
rect 563482 494161 563542 494221
rect 563602 494161 563662 494221
rect 563722 494161 563782 494221
rect 563842 494161 563902 494221
rect 563962 494161 564022 494221
rect 564082 494161 564142 494221
rect 564202 494161 564262 494221
rect 564322 494161 564382 494221
rect 564442 494161 564502 494221
rect 564562 494161 564622 494221
rect 564682 494161 564742 494221
rect 564802 494161 564862 494221
rect 564922 494161 564982 494221
rect 565042 494161 565102 494221
rect 565162 494161 565222 494221
rect 565282 494161 565342 494221
rect 565402 494161 565462 494221
rect 565522 494161 565582 494221
rect 565642 494161 565702 494221
rect 565762 494161 565822 494221
rect 565882 494161 565942 494221
rect 566002 494161 566062 494221
rect 566122 494161 566182 494221
rect 566242 494161 566302 494221
rect 566362 494161 566422 494221
rect 566482 494161 566542 494221
rect 566602 494161 566662 494221
rect 566722 494161 566782 494221
rect 566842 494161 566902 494221
rect 566962 494161 567022 494221
rect 567082 494161 567142 494221
rect 567202 494161 567262 494221
rect 567322 494161 567382 494221
rect 567442 494161 567502 494221
rect 567562 494161 567622 494221
rect 562102 494101 567622 494161
rect 562102 494041 562222 494101
rect 562282 494041 562342 494101
rect 562402 494041 562462 494101
rect 562522 494041 562582 494101
rect 562642 494041 562702 494101
rect 562762 494041 562822 494101
rect 562882 494041 562942 494101
rect 563002 494041 563062 494101
rect 563122 494041 563182 494101
rect 563242 494041 563302 494101
rect 563362 494041 563422 494101
rect 563482 494041 563542 494101
rect 563602 494041 563662 494101
rect 563722 494041 563782 494101
rect 563842 494041 563902 494101
rect 563962 494041 564022 494101
rect 564082 494041 564142 494101
rect 564202 494041 564262 494101
rect 564322 494041 564382 494101
rect 564442 494041 564502 494101
rect 564562 494041 564622 494101
rect 564682 494041 564742 494101
rect 564802 494041 564862 494101
rect 564922 494041 564982 494101
rect 565042 494041 565102 494101
rect 565162 494041 565222 494101
rect 565282 494041 565342 494101
rect 565402 494041 565462 494101
rect 565522 494041 565582 494101
rect 565642 494041 565702 494101
rect 565762 494041 565822 494101
rect 565882 494041 565942 494101
rect 566002 494041 566062 494101
rect 566122 494041 566182 494101
rect 566242 494041 566302 494101
rect 566362 494041 566422 494101
rect 566482 494041 566542 494101
rect 566602 494041 566662 494101
rect 566722 494041 566782 494101
rect 566842 494041 566902 494101
rect 566962 494041 567022 494101
rect 567082 494041 567142 494101
rect 567202 494041 567262 494101
rect 567322 494041 567382 494101
rect 567442 494041 567502 494101
rect 567562 494041 567622 494101
rect 562102 493981 567622 494041
rect 572272 494236 577792 494296
rect 572272 494176 572332 494236
rect 572392 494176 572452 494236
rect 572512 494176 572572 494236
rect 572632 494176 572692 494236
rect 572752 494176 572812 494236
rect 572872 494176 572932 494236
rect 572992 494176 573052 494236
rect 573112 494176 573172 494236
rect 573232 494176 573292 494236
rect 573352 494176 573412 494236
rect 573472 494176 573532 494236
rect 573592 494176 573652 494236
rect 573712 494176 573772 494236
rect 573832 494176 573892 494236
rect 573952 494176 574012 494236
rect 574072 494176 574132 494236
rect 574192 494176 574252 494236
rect 574312 494176 574372 494236
rect 574432 494176 574492 494236
rect 574552 494176 574612 494236
rect 574672 494176 574732 494236
rect 574792 494176 574852 494236
rect 574912 494176 574972 494236
rect 575032 494176 575092 494236
rect 575152 494176 575212 494236
rect 575272 494176 575332 494236
rect 575392 494176 575452 494236
rect 575512 494176 575572 494236
rect 575632 494176 575692 494236
rect 575752 494176 575812 494236
rect 575872 494176 575932 494236
rect 575992 494176 576052 494236
rect 576112 494176 576172 494236
rect 576232 494176 576292 494236
rect 576352 494176 576412 494236
rect 576472 494176 576532 494236
rect 576592 494176 576652 494236
rect 576712 494176 576772 494236
rect 576832 494176 576892 494236
rect 576952 494176 577012 494236
rect 577072 494176 577132 494236
rect 577192 494176 577252 494236
rect 577312 494176 577372 494236
rect 577432 494176 577492 494236
rect 577552 494176 577612 494236
rect 577672 494176 577792 494236
rect 572272 494116 577792 494176
rect 572272 494056 572332 494116
rect 572392 494056 572452 494116
rect 572512 494056 572572 494116
rect 572632 494056 572692 494116
rect 572752 494056 572812 494116
rect 572872 494056 572932 494116
rect 572992 494056 573052 494116
rect 573112 494056 573172 494116
rect 573232 494056 573292 494116
rect 573352 494056 573412 494116
rect 573472 494056 573532 494116
rect 573592 494056 573652 494116
rect 573712 494056 573772 494116
rect 573832 494056 573892 494116
rect 573952 494056 574012 494116
rect 574072 494056 574132 494116
rect 574192 494056 574252 494116
rect 574312 494056 574372 494116
rect 574432 494056 574492 494116
rect 574552 494056 574612 494116
rect 574672 494056 574732 494116
rect 574792 494056 574852 494116
rect 574912 494056 574972 494116
rect 575032 494056 575092 494116
rect 575152 494056 575212 494116
rect 575272 494056 575332 494116
rect 575392 494056 575452 494116
rect 575512 494056 575572 494116
rect 575632 494056 575692 494116
rect 575752 494056 575812 494116
rect 575872 494056 575932 494116
rect 575992 494056 576052 494116
rect 576112 494056 576172 494116
rect 576232 494056 576292 494116
rect 576352 494056 576412 494116
rect 576472 494056 576532 494116
rect 576592 494056 576652 494116
rect 576712 494056 576772 494116
rect 576832 494056 576892 494116
rect 576952 494056 577012 494116
rect 577072 494056 577132 494116
rect 577192 494056 577252 494116
rect 577312 494056 577372 494116
rect 577432 494056 577492 494116
rect 577552 494056 577612 494116
rect 577672 494056 577792 494116
rect 572272 493996 577792 494056
rect 562380 455440 567480 455520
rect 562380 455360 562480 455440
rect 562560 455360 562640 455440
rect 562720 455360 562800 455440
rect 562880 455360 562960 455440
rect 563040 455360 563120 455440
rect 563200 455360 563280 455440
rect 563360 455360 563440 455440
rect 563520 455360 563600 455440
rect 563680 455360 563760 455440
rect 563840 455360 563920 455440
rect 564000 455360 564080 455440
rect 564160 455360 564240 455440
rect 564320 455360 564400 455440
rect 564480 455360 564560 455440
rect 564640 455360 564720 455440
rect 564800 455360 564880 455440
rect 564960 455360 565040 455440
rect 565120 455360 565200 455440
rect 565280 455360 565360 455440
rect 565440 455360 565520 455440
rect 565600 455360 565680 455440
rect 565760 455360 565840 455440
rect 565920 455360 566000 455440
rect 566080 455360 566160 455440
rect 566240 455360 566320 455440
rect 566400 455360 566480 455440
rect 566560 455360 566640 455440
rect 566720 455360 566800 455440
rect 566880 455360 566960 455440
rect 567040 455360 567120 455440
rect 567200 455360 567280 455440
rect 567360 455360 567480 455440
rect 562380 455280 567480 455360
rect 562380 455200 562480 455280
rect 562560 455200 562640 455280
rect 562720 455200 562800 455280
rect 562880 455200 562960 455280
rect 563040 455200 563120 455280
rect 563200 455200 563280 455280
rect 563360 455200 563440 455280
rect 563520 455200 563600 455280
rect 563680 455200 563760 455280
rect 563840 455200 563920 455280
rect 564000 455200 564080 455280
rect 564160 455200 564240 455280
rect 564320 455200 564400 455280
rect 564480 455200 564560 455280
rect 564640 455200 564720 455280
rect 564800 455200 564880 455280
rect 564960 455200 565040 455280
rect 565120 455200 565200 455280
rect 565280 455200 565360 455280
rect 565440 455200 565520 455280
rect 565600 455200 565680 455280
rect 565760 455200 565840 455280
rect 565920 455200 566000 455280
rect 566080 455200 566160 455280
rect 566240 455200 566320 455280
rect 566400 455200 566480 455280
rect 566560 455200 566640 455280
rect 566720 455200 566800 455280
rect 566880 455200 566960 455280
rect 567040 455200 567120 455280
rect 567200 455200 567280 455280
rect 567360 455200 567480 455280
rect 562380 455160 567480 455200
rect 572540 455440 577640 455520
rect 572540 455360 572640 455440
rect 572720 455360 572800 455440
rect 572880 455360 572960 455440
rect 573040 455360 573120 455440
rect 573200 455360 573280 455440
rect 573360 455360 573440 455440
rect 573520 455360 573600 455440
rect 573680 455360 573760 455440
rect 573840 455360 573920 455440
rect 574000 455360 574080 455440
rect 574160 455360 574240 455440
rect 574320 455360 574400 455440
rect 574480 455360 574560 455440
rect 574640 455360 574720 455440
rect 574800 455360 574880 455440
rect 574960 455360 575040 455440
rect 575120 455360 575200 455440
rect 575280 455360 575360 455440
rect 575440 455360 575520 455440
rect 575600 455360 575680 455440
rect 575760 455360 575840 455440
rect 575920 455360 576000 455440
rect 576080 455360 576160 455440
rect 576240 455360 576320 455440
rect 576400 455360 576480 455440
rect 576560 455360 576640 455440
rect 576720 455360 576800 455440
rect 576880 455360 576960 455440
rect 577040 455360 577120 455440
rect 577200 455360 577280 455440
rect 577360 455360 577440 455440
rect 577520 455360 577640 455440
rect 572540 455280 577640 455360
rect 572540 455200 572640 455280
rect 572720 455200 572800 455280
rect 572880 455200 572960 455280
rect 573040 455200 573120 455280
rect 573200 455200 573280 455280
rect 573360 455200 573440 455280
rect 573520 455200 573600 455280
rect 573680 455200 573760 455280
rect 573840 455200 573920 455280
rect 574000 455200 574080 455280
rect 574160 455200 574240 455280
rect 574320 455200 574400 455280
rect 574480 455200 574560 455280
rect 574640 455200 574720 455280
rect 574800 455200 574880 455280
rect 574960 455200 575040 455280
rect 575120 455200 575200 455280
rect 575280 455200 575360 455280
rect 575440 455200 575520 455280
rect 575600 455200 575680 455280
rect 575760 455200 575840 455280
rect 575920 455200 576000 455280
rect 576080 455200 576160 455280
rect 576240 455200 576320 455280
rect 576400 455200 576480 455280
rect 576560 455200 576640 455280
rect 576720 455200 576800 455280
rect 576880 455200 576960 455280
rect 577040 455200 577120 455280
rect 577200 455200 577280 455280
rect 577360 455200 577440 455280
rect 577520 455200 577640 455280
rect 572540 455160 577640 455200
rect 562102 453919 567622 453979
rect 562102 453859 562222 453919
rect 562282 453859 562342 453919
rect 562402 453859 562462 453919
rect 562522 453859 562582 453919
rect 562642 453859 562702 453919
rect 562762 453859 562822 453919
rect 562882 453859 562942 453919
rect 563002 453859 563062 453919
rect 563122 453859 563182 453919
rect 563242 453859 563302 453919
rect 563362 453859 563422 453919
rect 563482 453859 563542 453919
rect 563602 453859 563662 453919
rect 563722 453859 563782 453919
rect 563842 453859 563902 453919
rect 563962 453859 564022 453919
rect 564082 453859 564142 453919
rect 564202 453859 564262 453919
rect 564322 453859 564382 453919
rect 564442 453859 564502 453919
rect 564562 453859 564622 453919
rect 564682 453859 564742 453919
rect 564802 453859 564862 453919
rect 564922 453859 564982 453919
rect 565042 453859 565102 453919
rect 565162 453859 565222 453919
rect 565282 453859 565342 453919
rect 565402 453859 565462 453919
rect 565522 453859 565582 453919
rect 565642 453859 565702 453919
rect 565762 453859 565822 453919
rect 565882 453859 565942 453919
rect 566002 453859 566062 453919
rect 566122 453859 566182 453919
rect 566242 453859 566302 453919
rect 566362 453859 566422 453919
rect 566482 453859 566542 453919
rect 566602 453859 566662 453919
rect 566722 453859 566782 453919
rect 566842 453859 566902 453919
rect 566962 453859 567022 453919
rect 567082 453859 567142 453919
rect 567202 453859 567262 453919
rect 567322 453859 567382 453919
rect 567442 453859 567502 453919
rect 567562 453859 567622 453919
rect 562102 453799 567622 453859
rect 562102 453739 562222 453799
rect 562282 453739 562342 453799
rect 562402 453739 562462 453799
rect 562522 453739 562582 453799
rect 562642 453739 562702 453799
rect 562762 453739 562822 453799
rect 562882 453739 562942 453799
rect 563002 453739 563062 453799
rect 563122 453739 563182 453799
rect 563242 453739 563302 453799
rect 563362 453739 563422 453799
rect 563482 453739 563542 453799
rect 563602 453739 563662 453799
rect 563722 453739 563782 453799
rect 563842 453739 563902 453799
rect 563962 453739 564022 453799
rect 564082 453739 564142 453799
rect 564202 453739 564262 453799
rect 564322 453739 564382 453799
rect 564442 453739 564502 453799
rect 564562 453739 564622 453799
rect 564682 453739 564742 453799
rect 564802 453739 564862 453799
rect 564922 453739 564982 453799
rect 565042 453739 565102 453799
rect 565162 453739 565222 453799
rect 565282 453739 565342 453799
rect 565402 453739 565462 453799
rect 565522 453739 565582 453799
rect 565642 453739 565702 453799
rect 565762 453739 565822 453799
rect 565882 453739 565942 453799
rect 566002 453739 566062 453799
rect 566122 453739 566182 453799
rect 566242 453739 566302 453799
rect 566362 453739 566422 453799
rect 566482 453739 566542 453799
rect 566602 453739 566662 453799
rect 566722 453739 566782 453799
rect 566842 453739 566902 453799
rect 566962 453739 567022 453799
rect 567082 453739 567142 453799
rect 567202 453739 567262 453799
rect 567322 453739 567382 453799
rect 567442 453739 567502 453799
rect 567562 453739 567622 453799
rect 562102 453679 567622 453739
rect 572272 453934 577792 453994
rect 572272 453874 572332 453934
rect 572392 453874 572452 453934
rect 572512 453874 572572 453934
rect 572632 453874 572692 453934
rect 572752 453874 572812 453934
rect 572872 453874 572932 453934
rect 572992 453874 573052 453934
rect 573112 453874 573172 453934
rect 573232 453874 573292 453934
rect 573352 453874 573412 453934
rect 573472 453874 573532 453934
rect 573592 453874 573652 453934
rect 573712 453874 573772 453934
rect 573832 453874 573892 453934
rect 573952 453874 574012 453934
rect 574072 453874 574132 453934
rect 574192 453874 574252 453934
rect 574312 453874 574372 453934
rect 574432 453874 574492 453934
rect 574552 453874 574612 453934
rect 574672 453874 574732 453934
rect 574792 453874 574852 453934
rect 574912 453874 574972 453934
rect 575032 453874 575092 453934
rect 575152 453874 575212 453934
rect 575272 453874 575332 453934
rect 575392 453874 575452 453934
rect 575512 453874 575572 453934
rect 575632 453874 575692 453934
rect 575752 453874 575812 453934
rect 575872 453874 575932 453934
rect 575992 453874 576052 453934
rect 576112 453874 576172 453934
rect 576232 453874 576292 453934
rect 576352 453874 576412 453934
rect 576472 453874 576532 453934
rect 576592 453874 576652 453934
rect 576712 453874 576772 453934
rect 576832 453874 576892 453934
rect 576952 453874 577012 453934
rect 577072 453874 577132 453934
rect 577192 453874 577252 453934
rect 577312 453874 577372 453934
rect 577432 453874 577492 453934
rect 577552 453874 577612 453934
rect 577672 453874 577792 453934
rect 572272 453814 577792 453874
rect 572272 453754 572332 453814
rect 572392 453754 572452 453814
rect 572512 453754 572572 453814
rect 572632 453754 572692 453814
rect 572752 453754 572812 453814
rect 572872 453754 572932 453814
rect 572992 453754 573052 453814
rect 573112 453754 573172 453814
rect 573232 453754 573292 453814
rect 573352 453754 573412 453814
rect 573472 453754 573532 453814
rect 573592 453754 573652 453814
rect 573712 453754 573772 453814
rect 573832 453754 573892 453814
rect 573952 453754 574012 453814
rect 574072 453754 574132 453814
rect 574192 453754 574252 453814
rect 574312 453754 574372 453814
rect 574432 453754 574492 453814
rect 574552 453754 574612 453814
rect 574672 453754 574732 453814
rect 574792 453754 574852 453814
rect 574912 453754 574972 453814
rect 575032 453754 575092 453814
rect 575152 453754 575212 453814
rect 575272 453754 575332 453814
rect 575392 453754 575452 453814
rect 575512 453754 575572 453814
rect 575632 453754 575692 453814
rect 575752 453754 575812 453814
rect 575872 453754 575932 453814
rect 575992 453754 576052 453814
rect 576112 453754 576172 453814
rect 576232 453754 576292 453814
rect 576352 453754 576412 453814
rect 576472 453754 576532 453814
rect 576592 453754 576652 453814
rect 576712 453754 576772 453814
rect 576832 453754 576892 453814
rect 576952 453754 577012 453814
rect 577072 453754 577132 453814
rect 577192 453754 577252 453814
rect 577312 453754 577372 453814
rect 577432 453754 577492 453814
rect 577552 453754 577612 453814
rect 577672 453754 577792 453814
rect 572272 453694 577792 453754
rect 524 -800 636 480
rect 1706 -800 1818 480
rect 2888 -800 3000 480
rect 4070 -800 4182 480
rect 5252 -800 5364 480
rect 6434 -800 6546 480
rect 7616 -800 7728 480
rect 8798 -800 8910 480
rect 9980 -800 10092 480
rect 11162 -800 11274 480
rect 12344 -800 12456 480
rect 13526 -800 13638 480
rect 14708 -800 14820 480
rect 15890 -800 16002 480
rect 17072 -800 17184 480
rect 18254 -800 18366 480
rect 19436 -800 19548 480
rect 20618 -800 20730 480
rect 21800 -800 21912 480
rect 22982 -800 23094 480
rect 24164 -800 24276 480
rect 25346 -800 25458 480
rect 26528 -800 26640 480
rect 27710 -800 27822 480
rect 28892 -800 29004 480
rect 30074 -800 30186 480
rect 31256 -800 31368 480
rect 32438 -800 32550 480
rect 33620 -800 33732 480
rect 34802 -800 34914 480
rect 35984 -800 36096 480
rect 37166 -800 37278 480
rect 38348 -800 38460 480
rect 39530 -800 39642 480
rect 40712 -800 40824 480
rect 41894 -800 42006 480
rect 43076 -800 43188 480
rect 44258 -800 44370 480
rect 45440 -800 45552 480
rect 46622 -800 46734 480
rect 47804 -800 47916 480
rect 48986 -800 49098 480
rect 50168 -800 50280 480
rect 51350 -800 51462 480
rect 52532 -800 52644 480
rect 53714 -800 53826 480
rect 54896 -800 55008 480
rect 56078 -800 56190 480
rect 57260 -800 57372 480
rect 58442 -800 58554 480
rect 59624 -800 59736 480
rect 60806 -800 60918 480
rect 61988 -800 62100 480
rect 63170 -800 63282 480
rect 64352 -800 64464 480
rect 65534 -800 65646 480
rect 66716 -800 66828 480
rect 67898 -800 68010 480
rect 69080 -800 69192 480
rect 70262 -800 70374 480
rect 71444 -800 71556 480
rect 72626 -800 72738 480
rect 73808 -800 73920 480
rect 74990 -800 75102 480
rect 76172 -800 76284 480
rect 77354 -800 77466 480
rect 78536 -800 78648 480
rect 79718 -800 79830 480
rect 80900 -800 81012 480
rect 82082 -800 82194 480
rect 83264 -800 83376 480
rect 84446 -800 84558 480
rect 85628 -800 85740 480
rect 86810 -800 86922 480
rect 87992 -800 88104 480
rect 89174 -800 89286 480
rect 90356 -800 90468 480
rect 91538 -800 91650 480
rect 92720 -800 92832 480
rect 93902 -800 94014 480
rect 95084 -800 95196 480
rect 96266 -800 96378 480
rect 97448 -800 97560 480
rect 98630 -800 98742 480
rect 99812 -800 99924 480
rect 100994 -800 101106 480
rect 102176 -800 102288 480
rect 103358 -800 103470 480
rect 104540 -800 104652 480
rect 105722 -800 105834 480
rect 106904 -800 107016 480
rect 108086 -800 108198 480
rect 109268 -800 109380 480
rect 110450 -800 110562 480
rect 111632 -800 111744 480
rect 112814 -800 112926 480
rect 113996 -800 114108 480
rect 115178 -800 115290 480
rect 116360 -800 116472 480
rect 117542 -800 117654 480
rect 118724 -800 118836 480
rect 119906 -800 120018 480
rect 121088 -800 121200 480
rect 122270 -800 122382 480
rect 123452 -800 123564 480
rect 124634 -800 124746 480
rect 125816 -800 125928 480
rect 126998 -800 127110 480
rect 128180 -800 128292 480
rect 129362 -800 129474 480
rect 130544 -800 130656 480
rect 131726 -800 131838 480
rect 132908 -800 133020 480
rect 134090 -800 134202 480
rect 135272 -800 135384 480
rect 136454 -800 136566 480
rect 137636 -800 137748 480
rect 138818 -800 138930 480
rect 140000 -800 140112 480
rect 141182 -800 141294 480
rect 142364 -800 142476 480
rect 143546 -800 143658 480
rect 144728 -800 144840 480
rect 145910 -800 146022 480
rect 147092 -800 147204 480
rect 148274 -800 148386 480
rect 149456 -800 149568 480
rect 150638 -800 150750 480
rect 151820 -800 151932 480
rect 153002 -800 153114 480
rect 154184 -800 154296 480
rect 155366 -800 155478 480
rect 156548 -800 156660 480
rect 157730 -800 157842 480
rect 158912 -800 159024 480
rect 160094 -800 160206 480
rect 161276 -800 161388 480
rect 162458 -800 162570 480
rect 163640 -800 163752 480
rect 164822 -800 164934 480
rect 166004 -800 166116 480
rect 167186 -800 167298 480
rect 168368 -800 168480 480
rect 169550 -800 169662 480
rect 170732 -800 170844 480
rect 171914 -800 172026 480
rect 173096 -800 173208 480
rect 174278 -800 174390 480
rect 175460 -800 175572 480
rect 176642 -800 176754 480
rect 177824 -800 177936 480
rect 179006 -800 179118 480
rect 180188 -800 180300 480
rect 181370 -800 181482 480
rect 182552 -800 182664 480
rect 183734 -800 183846 480
rect 184916 -800 185028 480
rect 186098 -800 186210 480
rect 187280 -800 187392 480
rect 188462 -800 188574 480
rect 189644 -800 189756 480
rect 190826 -800 190938 480
rect 192008 -800 192120 480
rect 193190 -800 193302 480
rect 194372 -800 194484 480
rect 195554 -800 195666 480
rect 196736 -800 196848 480
rect 197918 -800 198030 480
rect 199100 -800 199212 480
rect 200282 -800 200394 480
rect 201464 -800 201576 480
rect 202646 -800 202758 480
rect 203828 -800 203940 480
rect 205010 -800 205122 480
rect 206192 -800 206304 480
rect 207374 -800 207486 480
rect 208556 -800 208668 480
rect 209738 -800 209850 480
rect 210920 -800 211032 480
rect 212102 -800 212214 480
rect 213284 -800 213396 480
rect 214466 -800 214578 480
rect 215648 -800 215760 480
rect 216830 -800 216942 480
rect 218012 -800 218124 480
rect 219194 -800 219306 480
rect 220376 -800 220488 480
rect 221558 -800 221670 480
rect 222740 -800 222852 480
rect 223922 -800 224034 480
rect 225104 -800 225216 480
rect 226286 -800 226398 480
rect 227468 -800 227580 480
rect 228650 -800 228762 480
rect 229832 -800 229944 480
rect 231014 -800 231126 480
rect 232196 -800 232308 480
rect 233378 -800 233490 480
rect 234560 -800 234672 480
rect 235742 -800 235854 480
rect 236924 -800 237036 480
rect 238106 -800 238218 480
rect 239288 -800 239400 480
rect 240470 -800 240582 480
rect 241652 -800 241764 480
rect 242834 -800 242946 480
rect 244016 -800 244128 480
rect 245198 -800 245310 480
rect 246380 -800 246492 480
rect 247562 -800 247674 480
rect 248744 -800 248856 480
rect 249926 -800 250038 480
rect 251108 -800 251220 480
rect 252290 -800 252402 480
rect 253472 -800 253584 480
rect 254654 -800 254766 480
rect 255836 -800 255948 480
rect 257018 -800 257130 480
rect 258200 -800 258312 480
rect 259382 -800 259494 480
rect 260564 -800 260676 480
rect 261746 -800 261858 480
rect 262928 -800 263040 480
rect 264110 -800 264222 480
rect 265292 -800 265404 480
rect 266474 -800 266586 480
rect 267656 -800 267768 480
rect 268838 -800 268950 480
rect 270020 -800 270132 480
rect 271202 -800 271314 480
rect 272384 -800 272496 480
rect 273566 -800 273678 480
rect 274748 -800 274860 480
rect 275930 -800 276042 480
rect 277112 -800 277224 480
rect 278294 -800 278406 480
rect 279476 -800 279588 480
rect 280658 -800 280770 480
rect 281840 -800 281952 480
rect 283022 -800 283134 480
rect 284204 -800 284316 480
rect 285386 -800 285498 480
rect 286568 -800 286680 480
rect 287750 -800 287862 480
rect 288932 -800 289044 480
rect 290114 -800 290226 480
rect 291296 -800 291408 480
rect 292478 -800 292590 480
rect 293660 -800 293772 480
rect 294842 -800 294954 480
rect 296024 -800 296136 480
rect 297206 -800 297318 480
rect 298388 -800 298500 480
rect 299570 -800 299682 480
rect 300752 -800 300864 480
rect 301934 -800 302046 480
rect 303116 -800 303228 480
rect 304298 -800 304410 480
rect 305480 -800 305592 480
rect 306662 -800 306774 480
rect 307844 -800 307956 480
rect 309026 -800 309138 480
rect 310208 -800 310320 480
rect 311390 -800 311502 480
rect 312572 -800 312684 480
rect 313754 -800 313866 480
rect 314936 -800 315048 480
rect 316118 -800 316230 480
rect 317300 -800 317412 480
rect 318482 -800 318594 480
rect 319664 -800 319776 480
rect 320846 -800 320958 480
rect 322028 -800 322140 480
rect 323210 -800 323322 480
rect 324392 -800 324504 480
rect 325574 -800 325686 480
rect 326756 -800 326868 480
rect 327938 -800 328050 480
rect 329120 -800 329232 480
rect 330302 -800 330414 480
rect 331484 -800 331596 480
rect 332666 -800 332778 480
rect 333848 -800 333960 480
rect 335030 -800 335142 480
rect 336212 -800 336324 480
rect 337394 -800 337506 480
rect 338576 -800 338688 480
rect 339758 -800 339870 480
rect 340940 -800 341052 480
rect 342122 -800 342234 480
rect 343304 -800 343416 480
rect 344486 -800 344598 480
rect 345668 -800 345780 480
rect 346850 -800 346962 480
rect 348032 -800 348144 480
rect 349214 -800 349326 480
rect 350396 -800 350508 480
rect 351578 -800 351690 480
rect 352760 -800 352872 480
rect 353942 -800 354054 480
rect 355124 -800 355236 480
rect 356306 -800 356418 480
rect 357488 -800 357600 480
rect 358670 -800 358782 480
rect 359852 -800 359964 480
rect 361034 -800 361146 480
rect 362216 -800 362328 480
rect 363398 -800 363510 480
rect 364580 -800 364692 480
rect 365762 -800 365874 480
rect 366944 -800 367056 480
rect 368126 -800 368238 480
rect 369308 -800 369420 480
rect 370490 -800 370602 480
rect 371672 -800 371784 480
rect 372854 -800 372966 480
rect 374036 -800 374148 480
rect 375218 -800 375330 480
rect 376400 -800 376512 480
rect 377582 -800 377694 480
rect 378764 -800 378876 480
rect 379946 -800 380058 480
rect 381128 -800 381240 480
rect 382310 -800 382422 480
rect 383492 -800 383604 480
rect 384674 -800 384786 480
rect 385856 -800 385968 480
rect 387038 -800 387150 480
rect 388220 -800 388332 480
rect 389402 -800 389514 480
rect 390584 -800 390696 480
rect 391766 -800 391878 480
rect 392948 -800 393060 480
rect 394130 -800 394242 480
rect 395312 -800 395424 480
rect 396494 -800 396606 480
rect 397676 -800 397788 480
rect 398858 -800 398970 480
rect 400040 -800 400152 480
rect 401222 -800 401334 480
rect 402404 -800 402516 480
rect 403586 -800 403698 480
rect 404768 -800 404880 480
rect 405950 -800 406062 480
rect 407132 -800 407244 480
rect 408314 -800 408426 480
rect 409496 -800 409608 480
rect 410678 -800 410790 480
rect 411860 -800 411972 480
rect 413042 -800 413154 480
rect 414224 -800 414336 480
rect 415406 -800 415518 480
rect 416588 -800 416700 480
rect 417770 -800 417882 480
rect 418952 -800 419064 480
rect 420134 -800 420246 480
rect 421316 -800 421428 480
rect 422498 -800 422610 480
rect 423680 -800 423792 480
rect 424862 -800 424974 480
rect 426044 -800 426156 480
rect 427226 -800 427338 480
rect 428408 -800 428520 480
rect 429590 -800 429702 480
rect 430772 -800 430884 480
rect 431954 -800 432066 480
rect 433136 -800 433248 480
rect 434318 -800 434430 480
rect 435500 -800 435612 480
rect 436682 -800 436794 480
rect 437864 -800 437976 480
rect 439046 -800 439158 480
rect 440228 -800 440340 480
rect 441410 -800 441522 480
rect 442592 -800 442704 480
rect 443774 -800 443886 480
rect 444956 -800 445068 480
rect 446138 -800 446250 480
rect 447320 -800 447432 480
rect 448502 -800 448614 480
rect 449684 -800 449796 480
rect 450866 -800 450978 480
rect 452048 -800 452160 480
rect 453230 -800 453342 480
rect 454412 -800 454524 480
rect 455594 -800 455706 480
rect 456776 -800 456888 480
rect 457958 -800 458070 480
rect 459140 -800 459252 480
rect 460322 -800 460434 480
rect 461504 -800 461616 480
rect 462686 -800 462798 480
rect 463868 -800 463980 480
rect 465050 -800 465162 480
rect 466232 -800 466344 480
rect 467414 -800 467526 480
rect 468596 -800 468708 480
rect 469778 -800 469890 480
rect 470960 -800 471072 480
rect 472142 -800 472254 480
rect 473324 -800 473436 480
rect 474506 -800 474618 480
rect 475688 -800 475800 480
rect 476870 -800 476982 480
rect 478052 -800 478164 480
rect 479234 -800 479346 480
rect 480416 -800 480528 480
rect 481598 -800 481710 480
rect 482780 -800 482892 480
rect 483962 -800 484074 480
rect 485144 -800 485256 480
rect 486326 -800 486438 480
rect 487508 -800 487620 480
rect 488690 -800 488802 480
rect 489872 -800 489984 480
rect 491054 -800 491166 480
rect 492236 -800 492348 480
rect 493418 -800 493530 480
rect 494600 -800 494712 480
rect 495782 -800 495894 480
rect 496964 -800 497076 480
rect 498146 -800 498258 480
rect 499328 -800 499440 480
rect 500510 -800 500622 480
rect 501692 -800 501804 480
rect 502874 -800 502986 480
rect 504056 -800 504168 480
rect 505238 -800 505350 480
rect 506420 -800 506532 480
rect 507602 -800 507714 480
rect 508784 -800 508896 480
rect 509966 -800 510078 480
rect 511148 -800 511260 480
rect 512330 -800 512442 480
rect 513512 -800 513624 480
rect 514694 -800 514806 480
rect 515876 -800 515988 480
rect 517058 -800 517170 480
rect 518240 -800 518352 480
rect 519422 -800 519534 480
rect 520604 -800 520716 480
rect 521786 -800 521898 480
rect 522968 -800 523080 480
rect 524150 -800 524262 480
rect 525332 -800 525444 480
rect 526514 -800 526626 480
rect 527696 -800 527808 480
rect 528878 -800 528990 480
rect 530060 -800 530172 480
rect 531242 -800 531354 480
rect 532424 -800 532536 480
rect 533606 -800 533718 480
rect 534788 -800 534900 480
rect 535970 -800 536082 480
rect 537152 -800 537264 480
rect 538334 -800 538446 480
rect 539516 -800 539628 480
rect 540698 -800 540810 480
rect 541880 -800 541992 480
rect 543062 -800 543174 480
rect 544244 -800 544356 480
rect 545426 -800 545538 480
rect 546608 -800 546720 480
rect 547790 -800 547902 480
rect 548972 -800 549084 480
rect 550154 -800 550266 480
rect 551336 -800 551448 480
rect 552518 -800 552630 480
rect 553700 -800 553812 480
rect 554882 -800 554994 480
rect 556064 -800 556176 480
rect 557246 -800 557358 480
rect 558428 -800 558540 480
rect 559610 -800 559722 480
rect 560792 -800 560904 480
rect 561974 -800 562086 480
rect 563156 -800 563268 480
rect 564338 -800 564450 480
rect 565520 -800 565632 480
rect 566702 -800 566814 480
rect 567884 -800 567996 480
rect 569066 -800 569178 480
rect 570248 -800 570360 480
rect 571430 -800 571542 480
rect 572612 -800 572724 480
rect 573794 -800 573906 480
rect 574976 -800 575088 480
rect 576158 -800 576270 480
rect 577340 -800 577452 480
rect 578522 -800 578634 480
rect 579704 -800 579816 480
rect 580886 -800 580998 480
rect 582068 -800 582180 480
rect 583250 -800 583362 480
<< via2 >>
rect 562480 495662 562560 495742
rect 562640 495662 562720 495742
rect 562800 495662 562880 495742
rect 562960 495662 563040 495742
rect 563120 495662 563200 495742
rect 563280 495662 563360 495742
rect 563440 495662 563520 495742
rect 563600 495662 563680 495742
rect 563760 495662 563840 495742
rect 563920 495662 564000 495742
rect 564080 495662 564160 495742
rect 564240 495662 564320 495742
rect 564400 495662 564480 495742
rect 564560 495662 564640 495742
rect 564720 495662 564800 495742
rect 564880 495662 564960 495742
rect 565040 495662 565120 495742
rect 565200 495662 565280 495742
rect 565360 495662 565440 495742
rect 565520 495662 565600 495742
rect 565680 495662 565760 495742
rect 565840 495662 565920 495742
rect 566000 495662 566080 495742
rect 566160 495662 566240 495742
rect 566320 495662 566400 495742
rect 566480 495662 566560 495742
rect 566640 495662 566720 495742
rect 566800 495662 566880 495742
rect 566960 495662 567040 495742
rect 567120 495662 567200 495742
rect 567280 495662 567360 495742
rect 562480 495502 562560 495582
rect 562640 495502 562720 495582
rect 562800 495502 562880 495582
rect 562960 495502 563040 495582
rect 563120 495502 563200 495582
rect 563280 495502 563360 495582
rect 563440 495502 563520 495582
rect 563600 495502 563680 495582
rect 563760 495502 563840 495582
rect 563920 495502 564000 495582
rect 564080 495502 564160 495582
rect 564240 495502 564320 495582
rect 564400 495502 564480 495582
rect 564560 495502 564640 495582
rect 564720 495502 564800 495582
rect 564880 495502 564960 495582
rect 565040 495502 565120 495582
rect 565200 495502 565280 495582
rect 565360 495502 565440 495582
rect 565520 495502 565600 495582
rect 565680 495502 565760 495582
rect 565840 495502 565920 495582
rect 566000 495502 566080 495582
rect 566160 495502 566240 495582
rect 566320 495502 566400 495582
rect 566480 495502 566560 495582
rect 566640 495502 566720 495582
rect 566800 495502 566880 495582
rect 566960 495502 567040 495582
rect 567120 495502 567200 495582
rect 567280 495502 567360 495582
rect 572640 495662 572720 495742
rect 572800 495662 572880 495742
rect 572960 495662 573040 495742
rect 573120 495662 573200 495742
rect 573280 495662 573360 495742
rect 573440 495662 573520 495742
rect 573600 495662 573680 495742
rect 573760 495662 573840 495742
rect 573920 495662 574000 495742
rect 574080 495662 574160 495742
rect 574240 495662 574320 495742
rect 574400 495662 574480 495742
rect 574560 495662 574640 495742
rect 574720 495662 574800 495742
rect 574880 495662 574960 495742
rect 575040 495662 575120 495742
rect 575200 495662 575280 495742
rect 575360 495662 575440 495742
rect 575520 495662 575600 495742
rect 575680 495662 575760 495742
rect 575840 495662 575920 495742
rect 576000 495662 576080 495742
rect 576160 495662 576240 495742
rect 576320 495662 576400 495742
rect 576480 495662 576560 495742
rect 576640 495662 576720 495742
rect 576800 495662 576880 495742
rect 576960 495662 577040 495742
rect 577120 495662 577200 495742
rect 577280 495662 577360 495742
rect 577440 495662 577520 495742
rect 572640 495502 572720 495582
rect 572800 495502 572880 495582
rect 572960 495502 573040 495582
rect 573120 495502 573200 495582
rect 573280 495502 573360 495582
rect 573440 495502 573520 495582
rect 573600 495502 573680 495582
rect 573760 495502 573840 495582
rect 573920 495502 574000 495582
rect 574080 495502 574160 495582
rect 574240 495502 574320 495582
rect 574400 495502 574480 495582
rect 574560 495502 574640 495582
rect 574720 495502 574800 495582
rect 574880 495502 574960 495582
rect 575040 495502 575120 495582
rect 575200 495502 575280 495582
rect 575360 495502 575440 495582
rect 575520 495502 575600 495582
rect 575680 495502 575760 495582
rect 575840 495502 575920 495582
rect 576000 495502 576080 495582
rect 576160 495502 576240 495582
rect 576320 495502 576400 495582
rect 576480 495502 576560 495582
rect 576640 495502 576720 495582
rect 576800 495502 576880 495582
rect 576960 495502 577040 495582
rect 577120 495502 577200 495582
rect 577280 495502 577360 495582
rect 577440 495502 577520 495582
rect 562222 494161 562282 494221
rect 562342 494161 562402 494221
rect 562462 494161 562522 494221
rect 562582 494161 562642 494221
rect 562702 494161 562762 494221
rect 562822 494161 562882 494221
rect 562942 494161 563002 494221
rect 563062 494161 563122 494221
rect 563182 494161 563242 494221
rect 563302 494161 563362 494221
rect 563422 494161 563482 494221
rect 563542 494161 563602 494221
rect 563662 494161 563722 494221
rect 563782 494161 563842 494221
rect 563902 494161 563962 494221
rect 564022 494161 564082 494221
rect 564142 494161 564202 494221
rect 564262 494161 564322 494221
rect 564382 494161 564442 494221
rect 564502 494161 564562 494221
rect 564622 494161 564682 494221
rect 564742 494161 564802 494221
rect 564862 494161 564922 494221
rect 564982 494161 565042 494221
rect 565102 494161 565162 494221
rect 565222 494161 565282 494221
rect 565342 494161 565402 494221
rect 565462 494161 565522 494221
rect 565582 494161 565642 494221
rect 565702 494161 565762 494221
rect 565822 494161 565882 494221
rect 565942 494161 566002 494221
rect 566062 494161 566122 494221
rect 566182 494161 566242 494221
rect 566302 494161 566362 494221
rect 566422 494161 566482 494221
rect 566542 494161 566602 494221
rect 566662 494161 566722 494221
rect 566782 494161 566842 494221
rect 566902 494161 566962 494221
rect 567022 494161 567082 494221
rect 567142 494161 567202 494221
rect 567262 494161 567322 494221
rect 567382 494161 567442 494221
rect 567502 494161 567562 494221
rect 562222 494041 562282 494101
rect 562342 494041 562402 494101
rect 562462 494041 562522 494101
rect 562582 494041 562642 494101
rect 562702 494041 562762 494101
rect 562822 494041 562882 494101
rect 562942 494041 563002 494101
rect 563062 494041 563122 494101
rect 563182 494041 563242 494101
rect 563302 494041 563362 494101
rect 563422 494041 563482 494101
rect 563542 494041 563602 494101
rect 563662 494041 563722 494101
rect 563782 494041 563842 494101
rect 563902 494041 563962 494101
rect 564022 494041 564082 494101
rect 564142 494041 564202 494101
rect 564262 494041 564322 494101
rect 564382 494041 564442 494101
rect 564502 494041 564562 494101
rect 564622 494041 564682 494101
rect 564742 494041 564802 494101
rect 564862 494041 564922 494101
rect 564982 494041 565042 494101
rect 565102 494041 565162 494101
rect 565222 494041 565282 494101
rect 565342 494041 565402 494101
rect 565462 494041 565522 494101
rect 565582 494041 565642 494101
rect 565702 494041 565762 494101
rect 565822 494041 565882 494101
rect 565942 494041 566002 494101
rect 566062 494041 566122 494101
rect 566182 494041 566242 494101
rect 566302 494041 566362 494101
rect 566422 494041 566482 494101
rect 566542 494041 566602 494101
rect 566662 494041 566722 494101
rect 566782 494041 566842 494101
rect 566902 494041 566962 494101
rect 567022 494041 567082 494101
rect 567142 494041 567202 494101
rect 567262 494041 567322 494101
rect 567382 494041 567442 494101
rect 567502 494041 567562 494101
rect 572332 494176 572392 494236
rect 572452 494176 572512 494236
rect 572572 494176 572632 494236
rect 572692 494176 572752 494236
rect 572812 494176 572872 494236
rect 572932 494176 572992 494236
rect 573052 494176 573112 494236
rect 573172 494176 573232 494236
rect 573292 494176 573352 494236
rect 573412 494176 573472 494236
rect 573532 494176 573592 494236
rect 573652 494176 573712 494236
rect 573772 494176 573832 494236
rect 573892 494176 573952 494236
rect 574012 494176 574072 494236
rect 574132 494176 574192 494236
rect 574252 494176 574312 494236
rect 574372 494176 574432 494236
rect 574492 494176 574552 494236
rect 574612 494176 574672 494236
rect 574732 494176 574792 494236
rect 574852 494176 574912 494236
rect 574972 494176 575032 494236
rect 575092 494176 575152 494236
rect 575212 494176 575272 494236
rect 575332 494176 575392 494236
rect 575452 494176 575512 494236
rect 575572 494176 575632 494236
rect 575692 494176 575752 494236
rect 575812 494176 575872 494236
rect 575932 494176 575992 494236
rect 576052 494176 576112 494236
rect 576172 494176 576232 494236
rect 576292 494176 576352 494236
rect 576412 494176 576472 494236
rect 576532 494176 576592 494236
rect 576652 494176 576712 494236
rect 576772 494176 576832 494236
rect 576892 494176 576952 494236
rect 577012 494176 577072 494236
rect 577132 494176 577192 494236
rect 577252 494176 577312 494236
rect 577372 494176 577432 494236
rect 577492 494176 577552 494236
rect 577612 494176 577672 494236
rect 572332 494056 572392 494116
rect 572452 494056 572512 494116
rect 572572 494056 572632 494116
rect 572692 494056 572752 494116
rect 572812 494056 572872 494116
rect 572932 494056 572992 494116
rect 573052 494056 573112 494116
rect 573172 494056 573232 494116
rect 573292 494056 573352 494116
rect 573412 494056 573472 494116
rect 573532 494056 573592 494116
rect 573652 494056 573712 494116
rect 573772 494056 573832 494116
rect 573892 494056 573952 494116
rect 574012 494056 574072 494116
rect 574132 494056 574192 494116
rect 574252 494056 574312 494116
rect 574372 494056 574432 494116
rect 574492 494056 574552 494116
rect 574612 494056 574672 494116
rect 574732 494056 574792 494116
rect 574852 494056 574912 494116
rect 574972 494056 575032 494116
rect 575092 494056 575152 494116
rect 575212 494056 575272 494116
rect 575332 494056 575392 494116
rect 575452 494056 575512 494116
rect 575572 494056 575632 494116
rect 575692 494056 575752 494116
rect 575812 494056 575872 494116
rect 575932 494056 575992 494116
rect 576052 494056 576112 494116
rect 576172 494056 576232 494116
rect 576292 494056 576352 494116
rect 576412 494056 576472 494116
rect 576532 494056 576592 494116
rect 576652 494056 576712 494116
rect 576772 494056 576832 494116
rect 576892 494056 576952 494116
rect 577012 494056 577072 494116
rect 577132 494056 577192 494116
rect 577252 494056 577312 494116
rect 577372 494056 577432 494116
rect 577492 494056 577552 494116
rect 577612 494056 577672 494116
rect 562480 455360 562560 455440
rect 562640 455360 562720 455440
rect 562800 455360 562880 455440
rect 562960 455360 563040 455440
rect 563120 455360 563200 455440
rect 563280 455360 563360 455440
rect 563440 455360 563520 455440
rect 563600 455360 563680 455440
rect 563760 455360 563840 455440
rect 563920 455360 564000 455440
rect 564080 455360 564160 455440
rect 564240 455360 564320 455440
rect 564400 455360 564480 455440
rect 564560 455360 564640 455440
rect 564720 455360 564800 455440
rect 564880 455360 564960 455440
rect 565040 455360 565120 455440
rect 565200 455360 565280 455440
rect 565360 455360 565440 455440
rect 565520 455360 565600 455440
rect 565680 455360 565760 455440
rect 565840 455360 565920 455440
rect 566000 455360 566080 455440
rect 566160 455360 566240 455440
rect 566320 455360 566400 455440
rect 566480 455360 566560 455440
rect 566640 455360 566720 455440
rect 566800 455360 566880 455440
rect 566960 455360 567040 455440
rect 567120 455360 567200 455440
rect 567280 455360 567360 455440
rect 562480 455200 562560 455280
rect 562640 455200 562720 455280
rect 562800 455200 562880 455280
rect 562960 455200 563040 455280
rect 563120 455200 563200 455280
rect 563280 455200 563360 455280
rect 563440 455200 563520 455280
rect 563600 455200 563680 455280
rect 563760 455200 563840 455280
rect 563920 455200 564000 455280
rect 564080 455200 564160 455280
rect 564240 455200 564320 455280
rect 564400 455200 564480 455280
rect 564560 455200 564640 455280
rect 564720 455200 564800 455280
rect 564880 455200 564960 455280
rect 565040 455200 565120 455280
rect 565200 455200 565280 455280
rect 565360 455200 565440 455280
rect 565520 455200 565600 455280
rect 565680 455200 565760 455280
rect 565840 455200 565920 455280
rect 566000 455200 566080 455280
rect 566160 455200 566240 455280
rect 566320 455200 566400 455280
rect 566480 455200 566560 455280
rect 566640 455200 566720 455280
rect 566800 455200 566880 455280
rect 566960 455200 567040 455280
rect 567120 455200 567200 455280
rect 567280 455200 567360 455280
rect 572640 455360 572720 455440
rect 572800 455360 572880 455440
rect 572960 455360 573040 455440
rect 573120 455360 573200 455440
rect 573280 455360 573360 455440
rect 573440 455360 573520 455440
rect 573600 455360 573680 455440
rect 573760 455360 573840 455440
rect 573920 455360 574000 455440
rect 574080 455360 574160 455440
rect 574240 455360 574320 455440
rect 574400 455360 574480 455440
rect 574560 455360 574640 455440
rect 574720 455360 574800 455440
rect 574880 455360 574960 455440
rect 575040 455360 575120 455440
rect 575200 455360 575280 455440
rect 575360 455360 575440 455440
rect 575520 455360 575600 455440
rect 575680 455360 575760 455440
rect 575840 455360 575920 455440
rect 576000 455360 576080 455440
rect 576160 455360 576240 455440
rect 576320 455360 576400 455440
rect 576480 455360 576560 455440
rect 576640 455360 576720 455440
rect 576800 455360 576880 455440
rect 576960 455360 577040 455440
rect 577120 455360 577200 455440
rect 577280 455360 577360 455440
rect 577440 455360 577520 455440
rect 572640 455200 572720 455280
rect 572800 455200 572880 455280
rect 572960 455200 573040 455280
rect 573120 455200 573200 455280
rect 573280 455200 573360 455280
rect 573440 455200 573520 455280
rect 573600 455200 573680 455280
rect 573760 455200 573840 455280
rect 573920 455200 574000 455280
rect 574080 455200 574160 455280
rect 574240 455200 574320 455280
rect 574400 455200 574480 455280
rect 574560 455200 574640 455280
rect 574720 455200 574800 455280
rect 574880 455200 574960 455280
rect 575040 455200 575120 455280
rect 575200 455200 575280 455280
rect 575360 455200 575440 455280
rect 575520 455200 575600 455280
rect 575680 455200 575760 455280
rect 575840 455200 575920 455280
rect 576000 455200 576080 455280
rect 576160 455200 576240 455280
rect 576320 455200 576400 455280
rect 576480 455200 576560 455280
rect 576640 455200 576720 455280
rect 576800 455200 576880 455280
rect 576960 455200 577040 455280
rect 577120 455200 577200 455280
rect 577280 455200 577360 455280
rect 577440 455200 577520 455280
rect 562222 453859 562282 453919
rect 562342 453859 562402 453919
rect 562462 453859 562522 453919
rect 562582 453859 562642 453919
rect 562702 453859 562762 453919
rect 562822 453859 562882 453919
rect 562942 453859 563002 453919
rect 563062 453859 563122 453919
rect 563182 453859 563242 453919
rect 563302 453859 563362 453919
rect 563422 453859 563482 453919
rect 563542 453859 563602 453919
rect 563662 453859 563722 453919
rect 563782 453859 563842 453919
rect 563902 453859 563962 453919
rect 564022 453859 564082 453919
rect 564142 453859 564202 453919
rect 564262 453859 564322 453919
rect 564382 453859 564442 453919
rect 564502 453859 564562 453919
rect 564622 453859 564682 453919
rect 564742 453859 564802 453919
rect 564862 453859 564922 453919
rect 564982 453859 565042 453919
rect 565102 453859 565162 453919
rect 565222 453859 565282 453919
rect 565342 453859 565402 453919
rect 565462 453859 565522 453919
rect 565582 453859 565642 453919
rect 565702 453859 565762 453919
rect 565822 453859 565882 453919
rect 565942 453859 566002 453919
rect 566062 453859 566122 453919
rect 566182 453859 566242 453919
rect 566302 453859 566362 453919
rect 566422 453859 566482 453919
rect 566542 453859 566602 453919
rect 566662 453859 566722 453919
rect 566782 453859 566842 453919
rect 566902 453859 566962 453919
rect 567022 453859 567082 453919
rect 567142 453859 567202 453919
rect 567262 453859 567322 453919
rect 567382 453859 567442 453919
rect 567502 453859 567562 453919
rect 562222 453739 562282 453799
rect 562342 453739 562402 453799
rect 562462 453739 562522 453799
rect 562582 453739 562642 453799
rect 562702 453739 562762 453799
rect 562822 453739 562882 453799
rect 562942 453739 563002 453799
rect 563062 453739 563122 453799
rect 563182 453739 563242 453799
rect 563302 453739 563362 453799
rect 563422 453739 563482 453799
rect 563542 453739 563602 453799
rect 563662 453739 563722 453799
rect 563782 453739 563842 453799
rect 563902 453739 563962 453799
rect 564022 453739 564082 453799
rect 564142 453739 564202 453799
rect 564262 453739 564322 453799
rect 564382 453739 564442 453799
rect 564502 453739 564562 453799
rect 564622 453739 564682 453799
rect 564742 453739 564802 453799
rect 564862 453739 564922 453799
rect 564982 453739 565042 453799
rect 565102 453739 565162 453799
rect 565222 453739 565282 453799
rect 565342 453739 565402 453799
rect 565462 453739 565522 453799
rect 565582 453739 565642 453799
rect 565702 453739 565762 453799
rect 565822 453739 565882 453799
rect 565942 453739 566002 453799
rect 566062 453739 566122 453799
rect 566182 453739 566242 453799
rect 566302 453739 566362 453799
rect 566422 453739 566482 453799
rect 566542 453739 566602 453799
rect 566662 453739 566722 453799
rect 566782 453739 566842 453799
rect 566902 453739 566962 453799
rect 567022 453739 567082 453799
rect 567142 453739 567202 453799
rect 567262 453739 567322 453799
rect 567382 453739 567442 453799
rect 567502 453739 567562 453799
rect 572332 453874 572392 453934
rect 572452 453874 572512 453934
rect 572572 453874 572632 453934
rect 572692 453874 572752 453934
rect 572812 453874 572872 453934
rect 572932 453874 572992 453934
rect 573052 453874 573112 453934
rect 573172 453874 573232 453934
rect 573292 453874 573352 453934
rect 573412 453874 573472 453934
rect 573532 453874 573592 453934
rect 573652 453874 573712 453934
rect 573772 453874 573832 453934
rect 573892 453874 573952 453934
rect 574012 453874 574072 453934
rect 574132 453874 574192 453934
rect 574252 453874 574312 453934
rect 574372 453874 574432 453934
rect 574492 453874 574552 453934
rect 574612 453874 574672 453934
rect 574732 453874 574792 453934
rect 574852 453874 574912 453934
rect 574972 453874 575032 453934
rect 575092 453874 575152 453934
rect 575212 453874 575272 453934
rect 575332 453874 575392 453934
rect 575452 453874 575512 453934
rect 575572 453874 575632 453934
rect 575692 453874 575752 453934
rect 575812 453874 575872 453934
rect 575932 453874 575992 453934
rect 576052 453874 576112 453934
rect 576172 453874 576232 453934
rect 576292 453874 576352 453934
rect 576412 453874 576472 453934
rect 576532 453874 576592 453934
rect 576652 453874 576712 453934
rect 576772 453874 576832 453934
rect 576892 453874 576952 453934
rect 577012 453874 577072 453934
rect 577132 453874 577192 453934
rect 577252 453874 577312 453934
rect 577372 453874 577432 453934
rect 577492 453874 577552 453934
rect 577612 453874 577672 453934
rect 572332 453754 572392 453814
rect 572452 453754 572512 453814
rect 572572 453754 572632 453814
rect 572692 453754 572752 453814
rect 572812 453754 572872 453814
rect 572932 453754 572992 453814
rect 573052 453754 573112 453814
rect 573172 453754 573232 453814
rect 573292 453754 573352 453814
rect 573412 453754 573472 453814
rect 573532 453754 573592 453814
rect 573652 453754 573712 453814
rect 573772 453754 573832 453814
rect 573892 453754 573952 453814
rect 574012 453754 574072 453814
rect 574132 453754 574192 453814
rect 574252 453754 574312 453814
rect 574372 453754 574432 453814
rect 574492 453754 574552 453814
rect 574612 453754 574672 453814
rect 574732 453754 574792 453814
rect 574852 453754 574912 453814
rect 574972 453754 575032 453814
rect 575092 453754 575152 453814
rect 575212 453754 575272 453814
rect 575332 453754 575392 453814
rect 575452 453754 575512 453814
rect 575572 453754 575632 453814
rect 575692 453754 575752 453814
rect 575812 453754 575872 453814
rect 575932 453754 575992 453814
rect 576052 453754 576112 453814
rect 576172 453754 576232 453814
rect 576292 453754 576352 453814
rect 576412 453754 576472 453814
rect 576532 453754 576592 453814
rect 576652 453754 576712 453814
rect 576772 453754 576832 453814
rect 576892 453754 576952 453814
rect 577012 453754 577072 453814
rect 577132 453754 577192 453814
rect 577252 453754 577312 453814
rect 577372 453754 577432 453814
rect 577492 453754 577552 453814
rect 577612 453754 577672 453814
<< metal3 >>
rect 16194 702300 21194 704800
rect 68194 702300 73194 704800
rect 120194 702300 125194 704800
rect 165594 702300 170594 704800
rect 170894 697200 173094 704800
rect 170894 692600 171000 697200
rect 173000 692600 173094 697200
rect 170894 692300 173094 692600
rect 173394 697200 175594 704800
rect 175894 702300 180894 704800
rect 217294 702300 222294 704800
rect 173394 692600 173400 697200
rect 175400 692600 175594 697200
rect 173394 692300 175594 692600
rect 222594 697200 224794 704800
rect 222594 692600 222706 697200
rect 224706 692600 224794 697200
rect 222594 692300 224794 692600
rect 225094 697200 227294 704800
rect 227594 702300 232594 704800
rect 318994 702300 323994 704800
rect 225094 692600 225106 697200
rect 227106 692600 227294 697200
rect 225094 692300 227294 692600
rect 324294 697200 326494 704800
rect 324294 692600 324412 697200
rect 326412 692600 326494 697200
rect 324294 692300 326494 692600
rect 326794 697200 328994 704800
rect 329294 702300 334294 704800
rect 413394 702300 418394 704800
rect 465394 702400 470394 704800
rect 326794 692600 326812 697200
rect 328812 692600 328994 697200
rect 326794 692300 328994 692600
rect 510594 697360 515394 704800
rect 510594 692560 510654 697360
rect 515334 692560 515394 697360
rect 510594 692500 515394 692560
rect 520594 697360 525394 704800
rect 566594 697380 571594 704800
rect 520594 692560 520654 697360
rect 525334 692560 525394 697360
rect 520594 692500 525394 692560
rect -800 680242 1700 685242
rect 577380 677984 584800 682984
rect -800 643842 1660 648642
rect 562480 644524 584800 644584
rect 562480 639844 562600 644524
rect 567400 639844 584800 644524
rect 562480 639784 584800 639844
rect -800 633842 1660 638642
rect 562540 634524 584800 634584
rect 562540 629844 562600 634524
rect 567400 629844 584800 634524
rect 562540 629784 584800 629844
rect 583520 589472 584800 589584
rect 583520 588290 584800 588402
rect 583520 587108 584800 587220
rect 583520 585926 584800 586038
rect 583520 584744 584800 584856
rect 583520 583562 584800 583674
rect -800 559442 1660 564242
rect -800 549442 1660 554242
rect 582340 550562 584800 555362
rect 582340 540562 584800 545362
rect 477192 522892 483800 523098
rect 562388 522892 567660 523006
rect 477060 522862 567660 522892
rect 477060 522626 477192 522862
rect 477428 522626 477664 522862
rect 477900 522626 478136 522862
rect 478372 522626 478608 522862
rect 478844 522626 479080 522862
rect 479316 522626 479552 522862
rect 479788 522626 480024 522862
rect 480260 522626 480496 522862
rect 480732 522626 480968 522862
rect 481204 522626 481440 522862
rect 481676 522626 481912 522862
rect 482148 522626 482384 522862
rect 482620 522626 482856 522862
rect 483092 522626 483328 522862
rect 483564 522740 567660 522862
rect 483564 522626 562624 522740
rect 477060 522504 562624 522626
rect 562860 522504 563096 522740
rect 563332 522504 563568 522740
rect 563804 522504 564040 522740
rect 564276 522504 564512 522740
rect 564748 522504 564984 522740
rect 565220 522504 565456 522740
rect 565692 522504 565928 522740
rect 566164 522504 566400 522740
rect 566636 522504 566872 522740
rect 567108 522504 567660 522740
rect 477060 522390 567660 522504
rect 477060 522154 477192 522390
rect 477428 522154 477664 522390
rect 477900 522154 478136 522390
rect 478372 522154 478608 522390
rect 478844 522154 479080 522390
rect 479316 522154 479552 522390
rect 479788 522154 480024 522390
rect 480260 522154 480496 522390
rect 480732 522154 480968 522390
rect 481204 522154 481440 522390
rect 481676 522154 481912 522390
rect 482148 522154 482384 522390
rect 482620 522154 482856 522390
rect 483092 522154 483328 522390
rect 483564 522268 567660 522390
rect 483564 522154 562624 522268
rect 477060 522032 562624 522154
rect 562860 522032 563096 522268
rect 563332 522032 563568 522268
rect 563804 522032 564040 522268
rect 564276 522032 564512 522268
rect 564748 522032 564984 522268
rect 565220 522032 565456 522268
rect 565692 522032 565928 522268
rect 566164 522032 566400 522268
rect 566636 522032 566872 522268
rect 567108 522032 567660 522268
rect 477060 521918 567660 522032
rect 477060 521682 477192 521918
rect 477428 521682 477664 521918
rect 477900 521682 478136 521918
rect 478372 521682 478608 521918
rect 478844 521682 479080 521918
rect 479316 521682 479552 521918
rect 479788 521682 480024 521918
rect 480260 521682 480496 521918
rect 480732 521682 480968 521918
rect 481204 521682 481440 521918
rect 481676 521682 481912 521918
rect 482148 521682 482384 521918
rect 482620 521682 482856 521918
rect 483092 521682 483328 521918
rect 483564 521796 567660 521918
rect 483564 521682 562624 521796
rect 477060 521560 562624 521682
rect 562860 521560 563096 521796
rect 563332 521560 563568 521796
rect 563804 521560 564040 521796
rect 564276 521560 564512 521796
rect 564748 521560 564984 521796
rect 565220 521560 565456 521796
rect 565692 521560 565928 521796
rect 566164 521560 566400 521796
rect 566636 521560 566872 521796
rect 567108 521560 567660 521796
rect 477060 521446 567660 521560
rect 477060 521210 477192 521446
rect 477428 521210 477664 521446
rect 477900 521210 478136 521446
rect 478372 521210 478608 521446
rect 478844 521210 479080 521446
rect 479316 521210 479552 521446
rect 479788 521210 480024 521446
rect 480260 521210 480496 521446
rect 480732 521210 480968 521446
rect 481204 521210 481440 521446
rect 481676 521210 481912 521446
rect 482148 521210 482384 521446
rect 482620 521210 482856 521446
rect 483092 521210 483328 521446
rect 483564 521324 567660 521446
rect 483564 521210 562624 521324
rect 477060 521088 562624 521210
rect 562860 521088 563096 521324
rect 563332 521088 563568 521324
rect 563804 521088 564040 521324
rect 564276 521088 564512 521324
rect 564748 521088 564984 521324
rect 565220 521088 565456 521324
rect 565692 521088 565928 521324
rect 566164 521088 566400 521324
rect 566636 521088 566872 521324
rect 567108 521088 567660 521324
rect 477060 520974 567660 521088
rect 477060 520738 477192 520974
rect 477428 520738 477664 520974
rect 477900 520738 478136 520974
rect 478372 520738 478608 520974
rect 478844 520738 479080 520974
rect 479316 520738 479552 520974
rect 479788 520738 480024 520974
rect 480260 520738 480496 520974
rect 480732 520738 480968 520974
rect 481204 520738 481440 520974
rect 481676 520738 481912 520974
rect 482148 520738 482384 520974
rect 482620 520738 482856 520974
rect 483092 520738 483328 520974
rect 483564 520852 567660 520974
rect 483564 520738 562624 520852
rect 477060 520616 562624 520738
rect 562860 520616 563096 520852
rect 563332 520616 563568 520852
rect 563804 520616 564040 520852
rect 564276 520616 564512 520852
rect 564748 520616 564984 520852
rect 565220 520616 565456 520852
rect 565692 520616 565928 520852
rect 566164 520616 566400 520852
rect 566636 520616 566872 520852
rect 567108 520616 567660 520852
rect 477060 520502 567660 520616
rect 477060 520266 477192 520502
rect 477428 520266 477664 520502
rect 477900 520266 478136 520502
rect 478372 520266 478608 520502
rect 478844 520266 479080 520502
rect 479316 520266 479552 520502
rect 479788 520266 480024 520502
rect 480260 520266 480496 520502
rect 480732 520266 480968 520502
rect 481204 520266 481440 520502
rect 481676 520266 481912 520502
rect 482148 520266 482384 520502
rect 482620 520266 482856 520502
rect 483092 520266 483328 520502
rect 483564 520380 567660 520502
rect 483564 520266 562624 520380
rect 477060 520144 562624 520266
rect 562860 520144 563096 520380
rect 563332 520144 563568 520380
rect 563804 520144 564040 520380
rect 564276 520144 564512 520380
rect 564748 520144 564984 520380
rect 565220 520144 565456 520380
rect 565692 520144 565928 520380
rect 566164 520144 566400 520380
rect 566636 520144 566872 520380
rect 567108 520144 567660 520380
rect 477060 520030 567660 520144
rect 477060 519794 477192 520030
rect 477428 519794 477664 520030
rect 477900 519794 478136 520030
rect 478372 519794 478608 520030
rect 478844 519794 479080 520030
rect 479316 519794 479552 520030
rect 479788 519794 480024 520030
rect 480260 519794 480496 520030
rect 480732 519794 480968 520030
rect 481204 519794 481440 520030
rect 481676 519794 481912 520030
rect 482148 519794 482384 520030
rect 482620 519794 482856 520030
rect 483092 519794 483328 520030
rect 483564 519908 567660 520030
rect 483564 519794 562624 519908
rect 477060 519672 562624 519794
rect 562860 519672 563096 519908
rect 563332 519672 563568 519908
rect 563804 519672 564040 519908
rect 564276 519672 564512 519908
rect 564748 519672 564984 519908
rect 565220 519672 565456 519908
rect 565692 519672 565928 519908
rect 566164 519672 566400 519908
rect 566636 519672 566872 519908
rect 567108 519672 567660 519908
rect 477060 519558 567660 519672
rect 477060 519322 477192 519558
rect 477428 519322 477664 519558
rect 477900 519322 478136 519558
rect 478372 519322 478608 519558
rect 478844 519322 479080 519558
rect 479316 519322 479552 519558
rect 479788 519322 480024 519558
rect 480260 519322 480496 519558
rect 480732 519322 480968 519558
rect 481204 519322 481440 519558
rect 481676 519322 481912 519558
rect 482148 519322 482384 519558
rect 482620 519322 482856 519558
rect 483092 519322 483328 519558
rect 483564 519436 567660 519558
rect 483564 519322 562624 519436
rect 477060 519200 562624 519322
rect 562860 519200 563096 519436
rect 563332 519200 563568 519436
rect 563804 519200 564040 519436
rect 564276 519200 564512 519436
rect 564748 519200 564984 519436
rect 565220 519200 565456 519436
rect 565692 519200 565928 519436
rect 566164 519200 566400 519436
rect 566636 519200 566872 519436
rect 567108 519200 567660 519436
rect 477060 519086 567660 519200
rect 477060 518850 477192 519086
rect 477428 518850 477664 519086
rect 477900 518850 478136 519086
rect 478372 518850 478608 519086
rect 478844 518850 479080 519086
rect 479316 518850 479552 519086
rect 479788 518850 480024 519086
rect 480260 518850 480496 519086
rect 480732 518850 480968 519086
rect 481204 518850 481440 519086
rect 481676 518850 481912 519086
rect 482148 518850 482384 519086
rect 482620 518850 482856 519086
rect 483092 518850 483328 519086
rect 483564 518964 567660 519086
rect 483564 518850 562624 518964
rect 477060 518728 562624 518850
rect 562860 518728 563096 518964
rect 563332 518728 563568 518964
rect 563804 518728 564040 518964
rect 564276 518728 564512 518964
rect 564748 518728 564984 518964
rect 565220 518728 565456 518964
rect 565692 518728 565928 518964
rect 566164 518728 566400 518964
rect 566636 518728 566872 518964
rect 567108 518728 567660 518964
rect 477060 518614 567660 518728
rect 477060 518378 477192 518614
rect 477428 518378 477664 518614
rect 477900 518378 478136 518614
rect 478372 518378 478608 518614
rect 478844 518378 479080 518614
rect 479316 518378 479552 518614
rect 479788 518378 480024 518614
rect 480260 518378 480496 518614
rect 480732 518378 480968 518614
rect 481204 518378 481440 518614
rect 481676 518378 481912 518614
rect 482148 518378 482384 518614
rect 482620 518378 482856 518614
rect 483092 518378 483328 518614
rect 483564 518492 567660 518614
rect 483564 518378 562624 518492
rect 477060 518256 562624 518378
rect 562860 518256 563096 518492
rect 563332 518256 563568 518492
rect 563804 518256 564040 518492
rect 564276 518256 564512 518492
rect 564748 518256 564984 518492
rect 565220 518256 565456 518492
rect 565692 518256 565928 518492
rect 566164 518256 566400 518492
rect 566636 518256 566872 518492
rect 567108 518256 567660 518492
rect 477060 518142 567660 518256
rect 477060 517906 477192 518142
rect 477428 517906 477664 518142
rect 477900 517906 478136 518142
rect 478372 517906 478608 518142
rect 478844 517906 479080 518142
rect 479316 517906 479552 518142
rect 479788 517906 480024 518142
rect 480260 517906 480496 518142
rect 480732 517906 480968 518142
rect 481204 517906 481440 518142
rect 481676 517906 481912 518142
rect 482148 517906 482384 518142
rect 482620 517906 482856 518142
rect 483092 517906 483328 518142
rect 483564 518020 567660 518142
rect 483564 517906 562624 518020
rect 477060 517784 562624 517906
rect 562860 517784 563096 518020
rect 563332 517784 563568 518020
rect 563804 517784 564040 518020
rect 564276 517784 564512 518020
rect 564748 517784 564984 518020
rect 565220 517784 565456 518020
rect 565692 517784 565928 518020
rect 566164 517784 566400 518020
rect 566636 517784 566872 518020
rect 567108 517784 567660 518020
rect 477060 517670 567660 517784
rect 477060 517434 477192 517670
rect 477428 517434 477664 517670
rect 477900 517434 478136 517670
rect 478372 517434 478608 517670
rect 478844 517434 479080 517670
rect 479316 517434 479552 517670
rect 479788 517434 480024 517670
rect 480260 517434 480496 517670
rect 480732 517434 480968 517670
rect 481204 517434 481440 517670
rect 481676 517434 481912 517670
rect 482148 517434 482384 517670
rect 482620 517434 482856 517670
rect 483092 517434 483328 517670
rect 483564 517548 567660 517670
rect 483564 517434 562624 517548
rect 477060 517312 562624 517434
rect 562860 517312 563096 517548
rect 563332 517312 563568 517548
rect 563804 517312 564040 517548
rect 564276 517312 564512 517548
rect 564748 517312 564984 517548
rect 565220 517312 565456 517548
rect 565692 517312 565928 517548
rect 566164 517312 566400 517548
rect 566636 517312 566872 517548
rect 567108 517312 567660 517548
rect 477060 517198 567660 517312
rect 477060 516962 477192 517198
rect 477428 516962 477664 517198
rect 477900 516962 478136 517198
rect 478372 516962 478608 517198
rect 478844 516962 479080 517198
rect 479316 516962 479552 517198
rect 479788 516962 480024 517198
rect 480260 516962 480496 517198
rect 480732 516962 480968 517198
rect 481204 516962 481440 517198
rect 481676 516962 481912 517198
rect 482148 516962 482384 517198
rect 482620 516962 482856 517198
rect 483092 516962 483328 517198
rect 483564 517076 567660 517198
rect 483564 516962 562624 517076
rect 477060 516840 562624 516962
rect 562860 516840 563096 517076
rect 563332 516840 563568 517076
rect 563804 516840 564040 517076
rect 564276 516840 564512 517076
rect 564748 516840 564984 517076
rect 565220 516840 565456 517076
rect 565692 516840 565928 517076
rect 566164 516840 566400 517076
rect 566636 516840 566872 517076
rect 567108 516840 567660 517076
rect 477060 516726 567660 516840
rect 477060 516490 477192 516726
rect 477428 516490 477664 516726
rect 477900 516490 478136 516726
rect 478372 516490 478608 516726
rect 478844 516490 479080 516726
rect 479316 516490 479552 516726
rect 479788 516490 480024 516726
rect 480260 516490 480496 516726
rect 480732 516490 480968 516726
rect 481204 516490 481440 516726
rect 481676 516490 481912 516726
rect 482148 516490 482384 516726
rect 482620 516490 482856 516726
rect 483092 516490 483328 516726
rect 483564 516604 567660 516726
rect 483564 516490 562624 516604
rect 477060 516368 562624 516490
rect 562860 516368 563096 516604
rect 563332 516368 563568 516604
rect 563804 516368 564040 516604
rect 564276 516368 564512 516604
rect 564748 516368 564984 516604
rect 565220 516368 565456 516604
rect 565692 516368 565928 516604
rect 566164 516368 566400 516604
rect 566636 516368 566872 516604
rect 567108 516368 567660 516604
rect 477060 516226 567660 516368
rect -800 511530 480 511642
rect -800 510348 480 510460
rect -800 509166 480 509278
rect -800 507984 480 508096
rect -800 506802 480 506914
rect -800 505620 480 505732
rect 583520 500050 584800 500162
rect 583520 498868 584800 498980
rect 583520 497686 584800 497798
rect 583520 496504 584800 496616
rect 562380 495742 567480 495822
rect 562380 495662 562480 495742
rect 562560 495662 562640 495742
rect 562720 495662 562800 495742
rect 562880 495662 562960 495742
rect 563040 495662 563120 495742
rect 563200 495662 563280 495742
rect 563360 495662 563440 495742
rect 563520 495662 563600 495742
rect 563680 495662 563760 495742
rect 563840 495662 563920 495742
rect 564000 495662 564080 495742
rect 564160 495662 564240 495742
rect 564320 495662 564400 495742
rect 564480 495662 564560 495742
rect 564640 495662 564720 495742
rect 564800 495662 564880 495742
rect 564960 495662 565040 495742
rect 565120 495662 565200 495742
rect 565280 495662 565360 495742
rect 565440 495662 565520 495742
rect 565600 495662 565680 495742
rect 565760 495662 565840 495742
rect 565920 495662 566000 495742
rect 566080 495662 566160 495742
rect 566240 495662 566320 495742
rect 566400 495662 566480 495742
rect 566560 495662 566640 495742
rect 566720 495662 566800 495742
rect 566880 495662 566960 495742
rect 567040 495662 567120 495742
rect 567200 495662 567280 495742
rect 567360 495662 567480 495742
rect 562380 495582 567480 495662
rect 562380 495502 562480 495582
rect 562560 495502 562640 495582
rect 562720 495502 562800 495582
rect 562880 495502 562960 495582
rect 563040 495502 563120 495582
rect 563200 495502 563280 495582
rect 563360 495502 563440 495582
rect 563520 495502 563600 495582
rect 563680 495502 563760 495582
rect 563840 495502 563920 495582
rect 564000 495502 564080 495582
rect 564160 495502 564240 495582
rect 564320 495502 564400 495582
rect 564480 495502 564560 495582
rect 564640 495502 564720 495582
rect 564800 495502 564880 495582
rect 564960 495502 565040 495582
rect 565120 495502 565200 495582
rect 565280 495502 565360 495582
rect 565440 495502 565520 495582
rect 565600 495502 565680 495582
rect 565760 495502 565840 495582
rect 565920 495502 566000 495582
rect 566080 495502 566160 495582
rect 566240 495502 566320 495582
rect 566400 495502 566480 495582
rect 566560 495502 566640 495582
rect 566720 495502 566800 495582
rect 566880 495502 566960 495582
rect 567040 495502 567120 495582
rect 567200 495502 567280 495582
rect 567360 495502 567480 495582
rect 562380 495462 567480 495502
rect 572540 495742 577640 495822
rect 572540 495662 572640 495742
rect 572720 495662 572800 495742
rect 572880 495662 572960 495742
rect 573040 495662 573120 495742
rect 573200 495662 573280 495742
rect 573360 495662 573440 495742
rect 573520 495662 573600 495742
rect 573680 495662 573760 495742
rect 573840 495662 573920 495742
rect 574000 495662 574080 495742
rect 574160 495662 574240 495742
rect 574320 495662 574400 495742
rect 574480 495662 574560 495742
rect 574640 495662 574720 495742
rect 574800 495662 574880 495742
rect 574960 495662 575040 495742
rect 575120 495662 575200 495742
rect 575280 495662 575360 495742
rect 575440 495662 575520 495742
rect 575600 495662 575680 495742
rect 575760 495662 575840 495742
rect 575920 495662 576000 495742
rect 576080 495662 576160 495742
rect 576240 495662 576320 495742
rect 576400 495662 576480 495742
rect 576560 495662 576640 495742
rect 576720 495662 576800 495742
rect 576880 495662 576960 495742
rect 577040 495662 577120 495742
rect 577200 495662 577280 495742
rect 577360 495662 577440 495742
rect 577520 495662 577640 495742
rect 572540 495582 577640 495662
rect 572540 495502 572640 495582
rect 572720 495502 572800 495582
rect 572880 495502 572960 495582
rect 573040 495502 573120 495582
rect 573200 495502 573280 495582
rect 573360 495502 573440 495582
rect 573520 495502 573600 495582
rect 573680 495502 573760 495582
rect 573840 495502 573920 495582
rect 574000 495502 574080 495582
rect 574160 495502 574240 495582
rect 574320 495502 574400 495582
rect 574480 495502 574560 495582
rect 574640 495502 574720 495582
rect 574800 495502 574880 495582
rect 574960 495502 575040 495582
rect 575120 495502 575200 495582
rect 575280 495502 575360 495582
rect 575440 495502 575520 495582
rect 575600 495502 575680 495582
rect 575760 495502 575840 495582
rect 575920 495502 576000 495582
rect 576080 495502 576160 495582
rect 576240 495502 576320 495582
rect 576400 495502 576480 495582
rect 576560 495502 576640 495582
rect 576720 495502 576800 495582
rect 576880 495502 576960 495582
rect 577040 495502 577120 495582
rect 577200 495502 577280 495582
rect 577360 495502 577440 495582
rect 577520 495502 577640 495582
rect 572540 495462 577640 495502
rect 583520 495322 584800 495434
rect 511400 494528 583800 494600
rect 511400 494464 511616 494528
rect 511680 494464 511744 494528
rect 511808 494464 511872 494528
rect 511936 494464 512000 494528
rect 512064 494464 583800 494528
rect 511400 494400 583800 494464
rect 511400 494336 511616 494400
rect 511680 494336 511744 494400
rect 511808 494336 511872 494400
rect 511936 494336 512000 494400
rect 512064 494336 583800 494400
rect 511400 494272 583800 494336
rect 511400 494208 511616 494272
rect 511680 494208 511744 494272
rect 511808 494208 511872 494272
rect 511936 494208 512000 494272
rect 512064 494252 583800 494272
rect 512064 494236 584800 494252
rect 512064 494221 572332 494236
rect 512064 494208 562222 494221
rect 511400 494161 562222 494208
rect 562282 494161 562342 494221
rect 562402 494161 562462 494221
rect 562522 494161 562582 494221
rect 562642 494161 562702 494221
rect 562762 494161 562822 494221
rect 562882 494161 562942 494221
rect 563002 494161 563062 494221
rect 563122 494161 563182 494221
rect 563242 494161 563302 494221
rect 563362 494161 563422 494221
rect 563482 494161 563542 494221
rect 563602 494161 563662 494221
rect 563722 494161 563782 494221
rect 563842 494161 563902 494221
rect 563962 494161 564022 494221
rect 564082 494161 564142 494221
rect 564202 494161 564262 494221
rect 564322 494161 564382 494221
rect 564442 494161 564502 494221
rect 564562 494161 564622 494221
rect 564682 494161 564742 494221
rect 564802 494161 564862 494221
rect 564922 494161 564982 494221
rect 565042 494161 565102 494221
rect 565162 494161 565222 494221
rect 565282 494161 565342 494221
rect 565402 494161 565462 494221
rect 565522 494161 565582 494221
rect 565642 494161 565702 494221
rect 565762 494161 565822 494221
rect 565882 494161 565942 494221
rect 566002 494161 566062 494221
rect 566122 494161 566182 494221
rect 566242 494161 566302 494221
rect 566362 494161 566422 494221
rect 566482 494161 566542 494221
rect 566602 494161 566662 494221
rect 566722 494161 566782 494221
rect 566842 494161 566902 494221
rect 566962 494161 567022 494221
rect 567082 494161 567142 494221
rect 567202 494161 567262 494221
rect 567322 494161 567382 494221
rect 567442 494161 567502 494221
rect 567562 494176 572332 494221
rect 572392 494176 572452 494236
rect 572512 494176 572572 494236
rect 572632 494176 572692 494236
rect 572752 494176 572812 494236
rect 572872 494176 572932 494236
rect 572992 494176 573052 494236
rect 573112 494176 573172 494236
rect 573232 494176 573292 494236
rect 573352 494176 573412 494236
rect 573472 494176 573532 494236
rect 573592 494176 573652 494236
rect 573712 494176 573772 494236
rect 573832 494176 573892 494236
rect 573952 494176 574012 494236
rect 574072 494176 574132 494236
rect 574192 494176 574252 494236
rect 574312 494176 574372 494236
rect 574432 494176 574492 494236
rect 574552 494176 574612 494236
rect 574672 494176 574732 494236
rect 574792 494176 574852 494236
rect 574912 494176 574972 494236
rect 575032 494176 575092 494236
rect 575152 494176 575212 494236
rect 575272 494176 575332 494236
rect 575392 494176 575452 494236
rect 575512 494176 575572 494236
rect 575632 494176 575692 494236
rect 575752 494176 575812 494236
rect 575872 494176 575932 494236
rect 575992 494176 576052 494236
rect 576112 494176 576172 494236
rect 576232 494176 576292 494236
rect 576352 494176 576412 494236
rect 576472 494176 576532 494236
rect 576592 494176 576652 494236
rect 576712 494176 576772 494236
rect 576832 494176 576892 494236
rect 576952 494176 577012 494236
rect 577072 494176 577132 494236
rect 577192 494176 577252 494236
rect 577312 494176 577372 494236
rect 577432 494176 577492 494236
rect 577552 494176 577612 494236
rect 577672 494176 584800 494236
rect 567562 494161 584800 494176
rect 511400 494144 584800 494161
rect 511400 494080 511616 494144
rect 511680 494080 511744 494144
rect 511808 494080 511872 494144
rect 511936 494080 512000 494144
rect 512064 494140 584800 494144
rect 512064 494116 583800 494140
rect 512064 494101 572332 494116
rect 512064 494080 562222 494101
rect 511400 494041 562222 494080
rect 562282 494041 562342 494101
rect 562402 494041 562462 494101
rect 562522 494041 562582 494101
rect 562642 494041 562702 494101
rect 562762 494041 562822 494101
rect 562882 494041 562942 494101
rect 563002 494041 563062 494101
rect 563122 494041 563182 494101
rect 563242 494041 563302 494101
rect 563362 494041 563422 494101
rect 563482 494041 563542 494101
rect 563602 494041 563662 494101
rect 563722 494041 563782 494101
rect 563842 494041 563902 494101
rect 563962 494041 564022 494101
rect 564082 494041 564142 494101
rect 564202 494041 564262 494101
rect 564322 494041 564382 494101
rect 564442 494041 564502 494101
rect 564562 494041 564622 494101
rect 564682 494041 564742 494101
rect 564802 494041 564862 494101
rect 564922 494041 564982 494101
rect 565042 494041 565102 494101
rect 565162 494041 565222 494101
rect 565282 494041 565342 494101
rect 565402 494041 565462 494101
rect 565522 494041 565582 494101
rect 565642 494041 565702 494101
rect 565762 494041 565822 494101
rect 565882 494041 565942 494101
rect 566002 494041 566062 494101
rect 566122 494041 566182 494101
rect 566242 494041 566302 494101
rect 566362 494041 566422 494101
rect 566482 494041 566542 494101
rect 566602 494041 566662 494101
rect 566722 494041 566782 494101
rect 566842 494041 566902 494101
rect 566962 494041 567022 494101
rect 567082 494041 567142 494101
rect 567202 494041 567262 494101
rect 567322 494041 567382 494101
rect 567442 494041 567502 494101
rect 567562 494056 572332 494101
rect 572392 494056 572452 494116
rect 572512 494056 572572 494116
rect 572632 494056 572692 494116
rect 572752 494056 572812 494116
rect 572872 494056 572932 494116
rect 572992 494056 573052 494116
rect 573112 494056 573172 494116
rect 573232 494056 573292 494116
rect 573352 494056 573412 494116
rect 573472 494056 573532 494116
rect 573592 494056 573652 494116
rect 573712 494056 573772 494116
rect 573832 494056 573892 494116
rect 573952 494056 574012 494116
rect 574072 494056 574132 494116
rect 574192 494056 574252 494116
rect 574312 494056 574372 494116
rect 574432 494056 574492 494116
rect 574552 494056 574612 494116
rect 574672 494056 574732 494116
rect 574792 494056 574852 494116
rect 574912 494056 574972 494116
rect 575032 494056 575092 494116
rect 575152 494056 575212 494116
rect 575272 494056 575332 494116
rect 575392 494056 575452 494116
rect 575512 494056 575572 494116
rect 575632 494056 575692 494116
rect 575752 494056 575812 494116
rect 575872 494056 575932 494116
rect 575992 494056 576052 494116
rect 576112 494056 576172 494116
rect 576232 494056 576292 494116
rect 576352 494056 576412 494116
rect 576472 494056 576532 494116
rect 576592 494056 576652 494116
rect 576712 494056 576772 494116
rect 576832 494056 576892 494116
rect 576952 494056 577012 494116
rect 577072 494056 577132 494116
rect 577192 494056 577252 494116
rect 577312 494056 577372 494116
rect 577432 494056 577492 494116
rect 577552 494056 577612 494116
rect 577672 494056 583800 494116
rect 567562 494041 583800 494056
rect 511400 494016 583800 494041
rect 511400 493952 511616 494016
rect 511680 493952 511744 494016
rect 511808 493952 511872 494016
rect 511936 493952 512000 494016
rect 512064 493952 583800 494016
rect 511400 493888 583800 493952
rect 511400 493824 511616 493888
rect 511680 493824 511744 493888
rect 511808 493824 511872 493888
rect 511936 493824 512000 493888
rect 512064 493824 583800 493888
rect 511400 493800 583800 493824
rect 572536 484236 577492 484272
rect 536504 483800 578504 484236
rect 536504 483564 572772 483800
rect 573008 483564 573244 483800
rect 573480 483564 573716 483800
rect 573952 483564 574188 483800
rect 574424 483564 574660 483800
rect 574896 483564 575132 483800
rect 575368 483564 575604 483800
rect 575840 483564 576076 483800
rect 576312 483564 576548 483800
rect 576784 483564 577020 483800
rect 577256 483564 578504 483800
rect 536504 483328 578504 483564
rect 536504 483092 572772 483328
rect 573008 483092 573244 483328
rect 573480 483092 573716 483328
rect 573952 483092 574188 483328
rect 574424 483092 574660 483328
rect 574896 483092 575132 483328
rect 575368 483092 575604 483328
rect 575840 483092 576076 483328
rect 576312 483092 576548 483328
rect 576784 483092 577020 483328
rect 577256 483092 578504 483328
rect 536504 482856 578504 483092
rect 536504 482620 572772 482856
rect 573008 482620 573244 482856
rect 573480 482620 573716 482856
rect 573952 482620 574188 482856
rect 574424 482620 574660 482856
rect 574896 482620 575132 482856
rect 575368 482620 575604 482856
rect 575840 482620 576076 482856
rect 576312 482620 576548 482856
rect 576784 482620 577020 482856
rect 577256 482620 578504 482856
rect 536504 482384 578504 482620
rect 536504 482148 572772 482384
rect 573008 482148 573244 482384
rect 573480 482148 573716 482384
rect 573952 482148 574188 482384
rect 574424 482148 574660 482384
rect 574896 482148 575132 482384
rect 575368 482148 575604 482384
rect 575840 482148 576076 482384
rect 576312 482148 576548 482384
rect 576784 482148 577020 482384
rect 577256 482148 578504 482384
rect 536504 481912 578504 482148
rect 536504 481676 572772 481912
rect 573008 481676 573244 481912
rect 573480 481676 573716 481912
rect 573952 481676 574188 481912
rect 574424 481676 574660 481912
rect 574896 481676 575132 481912
rect 575368 481676 575604 481912
rect 575840 481676 576076 481912
rect 576312 481676 576548 481912
rect 576784 481676 577020 481912
rect 577256 481676 578504 481912
rect 536504 481440 578504 481676
rect 536504 481204 572772 481440
rect 573008 481204 573244 481440
rect 573480 481204 573716 481440
rect 573952 481204 574188 481440
rect 574424 481204 574660 481440
rect 574896 481204 575132 481440
rect 575368 481204 575604 481440
rect 575840 481204 576076 481440
rect 576312 481204 576548 481440
rect 576784 481204 577020 481440
rect 577256 481204 578504 481440
rect 536504 480968 578504 481204
rect 536504 480732 572772 480968
rect 573008 480732 573244 480968
rect 573480 480732 573716 480968
rect 573952 480732 574188 480968
rect 574424 480732 574660 480968
rect 574896 480732 575132 480968
rect 575368 480732 575604 480968
rect 575840 480732 576076 480968
rect 576312 480732 576548 480968
rect 576784 480732 577020 480968
rect 577256 480732 578504 480968
rect 536504 480496 578504 480732
rect 536504 480260 572772 480496
rect 573008 480260 573244 480496
rect 573480 480260 573716 480496
rect 573952 480260 574188 480496
rect 574424 480260 574660 480496
rect 574896 480260 575132 480496
rect 575368 480260 575604 480496
rect 575840 480260 576076 480496
rect 576312 480260 576548 480496
rect 576784 480260 577020 480496
rect 577256 480260 578504 480496
rect 536504 480024 578504 480260
rect 536504 479788 572772 480024
rect 573008 479788 573244 480024
rect 573480 479788 573716 480024
rect 573952 479788 574188 480024
rect 574424 479788 574660 480024
rect 574896 479788 575132 480024
rect 575368 479788 575604 480024
rect 575840 479788 576076 480024
rect 576312 479788 576548 480024
rect 576784 479788 577020 480024
rect 577256 479788 578504 480024
rect 536504 479552 578504 479788
rect 536504 479316 572772 479552
rect 573008 479316 573244 479552
rect 573480 479316 573716 479552
rect 573952 479316 574188 479552
rect 574424 479316 574660 479552
rect 574896 479316 575132 479552
rect 575368 479316 575604 479552
rect 575840 479316 576076 479552
rect 576312 479316 576548 479552
rect 576784 479316 577020 479552
rect 577256 479316 578504 479552
rect 536504 479080 578504 479316
rect 536504 478844 572772 479080
rect 573008 478844 573244 479080
rect 573480 478844 573716 479080
rect 573952 478844 574188 479080
rect 574424 478844 574660 479080
rect 574896 478844 575132 479080
rect 575368 478844 575604 479080
rect 575840 478844 576076 479080
rect 576312 478844 576548 479080
rect 576784 478844 577020 479080
rect 577256 478844 578504 479080
rect 536504 478608 578504 478844
rect 536504 478372 572772 478608
rect 573008 478372 573244 478608
rect 573480 478372 573716 478608
rect 573952 478372 574188 478608
rect 574424 478372 574660 478608
rect 574896 478372 575132 478608
rect 575368 478372 575604 478608
rect 575840 478372 576076 478608
rect 576312 478372 576548 478608
rect 576784 478372 577020 478608
rect 577256 478372 578504 478608
rect 536504 478136 578504 478372
rect 536504 477900 572772 478136
rect 573008 477900 573244 478136
rect 573480 477900 573716 478136
rect 573952 477900 574188 478136
rect 574424 477900 574660 478136
rect 574896 477900 575132 478136
rect 575368 477900 575604 478136
rect 575840 477900 576076 478136
rect 576312 477900 576548 478136
rect 576784 477900 577020 478136
rect 577256 477900 578504 478136
rect 536504 477580 578504 477900
rect -800 468308 480 468420
rect -800 467126 480 467238
rect -800 465944 480 466056
rect -800 464762 480 464874
rect -800 463580 480 463692
rect -800 462398 480 462510
rect 583520 455628 584800 455740
rect 562380 455440 567480 455520
rect 562380 455360 562480 455440
rect 562560 455360 562640 455440
rect 562720 455360 562800 455440
rect 562880 455360 562960 455440
rect 563040 455360 563120 455440
rect 563200 455360 563280 455440
rect 563360 455360 563440 455440
rect 563520 455360 563600 455440
rect 563680 455360 563760 455440
rect 563840 455360 563920 455440
rect 564000 455360 564080 455440
rect 564160 455360 564240 455440
rect 564320 455360 564400 455440
rect 564480 455360 564560 455440
rect 564640 455360 564720 455440
rect 564800 455360 564880 455440
rect 564960 455360 565040 455440
rect 565120 455360 565200 455440
rect 565280 455360 565360 455440
rect 565440 455360 565520 455440
rect 565600 455360 565680 455440
rect 565760 455360 565840 455440
rect 565920 455360 566000 455440
rect 566080 455360 566160 455440
rect 566240 455360 566320 455440
rect 566400 455360 566480 455440
rect 566560 455360 566640 455440
rect 566720 455360 566800 455440
rect 566880 455360 566960 455440
rect 567040 455360 567120 455440
rect 567200 455360 567280 455440
rect 567360 455360 567480 455440
rect 562380 455280 567480 455360
rect 562380 455200 562480 455280
rect 562560 455200 562640 455280
rect 562720 455200 562800 455280
rect 562880 455200 562960 455280
rect 563040 455200 563120 455280
rect 563200 455200 563280 455280
rect 563360 455200 563440 455280
rect 563520 455200 563600 455280
rect 563680 455200 563760 455280
rect 563840 455200 563920 455280
rect 564000 455200 564080 455280
rect 564160 455200 564240 455280
rect 564320 455200 564400 455280
rect 564480 455200 564560 455280
rect 564640 455200 564720 455280
rect 564800 455200 564880 455280
rect 564960 455200 565040 455280
rect 565120 455200 565200 455280
rect 565280 455200 565360 455280
rect 565440 455200 565520 455280
rect 565600 455200 565680 455280
rect 565760 455200 565840 455280
rect 565920 455200 566000 455280
rect 566080 455200 566160 455280
rect 566240 455200 566320 455280
rect 566400 455200 566480 455280
rect 566560 455200 566640 455280
rect 566720 455200 566800 455280
rect 566880 455200 566960 455280
rect 567040 455200 567120 455280
rect 567200 455200 567280 455280
rect 567360 455200 567480 455280
rect 562380 455160 567480 455200
rect 572540 455440 577640 455520
rect 572540 455360 572640 455440
rect 572720 455360 572800 455440
rect 572880 455360 572960 455440
rect 573040 455360 573120 455440
rect 573200 455360 573280 455440
rect 573360 455360 573440 455440
rect 573520 455360 573600 455440
rect 573680 455360 573760 455440
rect 573840 455360 573920 455440
rect 574000 455360 574080 455440
rect 574160 455360 574240 455440
rect 574320 455360 574400 455440
rect 574480 455360 574560 455440
rect 574640 455360 574720 455440
rect 574800 455360 574880 455440
rect 574960 455360 575040 455440
rect 575120 455360 575200 455440
rect 575280 455360 575360 455440
rect 575440 455360 575520 455440
rect 575600 455360 575680 455440
rect 575760 455360 575840 455440
rect 575920 455360 576000 455440
rect 576080 455360 576160 455440
rect 576240 455360 576320 455440
rect 576400 455360 576480 455440
rect 576560 455360 576640 455440
rect 576720 455360 576800 455440
rect 576880 455360 576960 455440
rect 577040 455360 577120 455440
rect 577200 455360 577280 455440
rect 577360 455360 577440 455440
rect 577520 455360 577640 455440
rect 572540 455280 577640 455360
rect 572540 455200 572640 455280
rect 572720 455200 572800 455280
rect 572880 455200 572960 455280
rect 573040 455200 573120 455280
rect 573200 455200 573280 455280
rect 573360 455200 573440 455280
rect 573520 455200 573600 455280
rect 573680 455200 573760 455280
rect 573840 455200 573920 455280
rect 574000 455200 574080 455280
rect 574160 455200 574240 455280
rect 574320 455200 574400 455280
rect 574480 455200 574560 455280
rect 574640 455200 574720 455280
rect 574800 455200 574880 455280
rect 574960 455200 575040 455280
rect 575120 455200 575200 455280
rect 575280 455200 575360 455280
rect 575440 455200 575520 455280
rect 575600 455200 575680 455280
rect 575760 455200 575840 455280
rect 575920 455200 576000 455280
rect 576080 455200 576160 455280
rect 576240 455200 576320 455280
rect 576400 455200 576480 455280
rect 576560 455200 576640 455280
rect 576720 455200 576800 455280
rect 576880 455200 576960 455280
rect 577040 455200 577120 455280
rect 577200 455200 577280 455280
rect 577360 455200 577440 455280
rect 577520 455200 577640 455280
rect 572540 455160 577640 455200
rect 583520 454446 584800 454558
rect 514788 453934 582788 454156
rect 514788 453919 572332 453934
rect 514788 453859 562222 453919
rect 562282 453859 562342 453919
rect 562402 453859 562462 453919
rect 562522 453859 562582 453919
rect 562642 453859 562702 453919
rect 562762 453859 562822 453919
rect 562882 453859 562942 453919
rect 563002 453859 563062 453919
rect 563122 453859 563182 453919
rect 563242 453859 563302 453919
rect 563362 453859 563422 453919
rect 563482 453859 563542 453919
rect 563602 453859 563662 453919
rect 563722 453859 563782 453919
rect 563842 453859 563902 453919
rect 563962 453859 564022 453919
rect 564082 453859 564142 453919
rect 564202 453859 564262 453919
rect 564322 453859 564382 453919
rect 564442 453859 564502 453919
rect 564562 453859 564622 453919
rect 564682 453859 564742 453919
rect 564802 453859 564862 453919
rect 564922 453859 564982 453919
rect 565042 453859 565102 453919
rect 565162 453859 565222 453919
rect 565282 453859 565342 453919
rect 565402 453859 565462 453919
rect 565522 453859 565582 453919
rect 565642 453859 565702 453919
rect 565762 453859 565822 453919
rect 565882 453859 565942 453919
rect 566002 453859 566062 453919
rect 566122 453859 566182 453919
rect 566242 453859 566302 453919
rect 566362 453859 566422 453919
rect 566482 453859 566542 453919
rect 566602 453859 566662 453919
rect 566722 453859 566782 453919
rect 566842 453859 566902 453919
rect 566962 453859 567022 453919
rect 567082 453859 567142 453919
rect 567202 453859 567262 453919
rect 567322 453859 567382 453919
rect 567442 453859 567502 453919
rect 567562 453874 572332 453919
rect 572392 453874 572452 453934
rect 572512 453874 572572 453934
rect 572632 453874 572692 453934
rect 572752 453874 572812 453934
rect 572872 453874 572932 453934
rect 572992 453874 573052 453934
rect 573112 453874 573172 453934
rect 573232 453874 573292 453934
rect 573352 453874 573412 453934
rect 573472 453874 573532 453934
rect 573592 453874 573652 453934
rect 573712 453874 573772 453934
rect 573832 453874 573892 453934
rect 573952 453874 574012 453934
rect 574072 453874 574132 453934
rect 574192 453874 574252 453934
rect 574312 453874 574372 453934
rect 574432 453874 574492 453934
rect 574552 453874 574612 453934
rect 574672 453874 574732 453934
rect 574792 453874 574852 453934
rect 574912 453874 574972 453934
rect 575032 453874 575092 453934
rect 575152 453874 575212 453934
rect 575272 453874 575332 453934
rect 575392 453874 575452 453934
rect 575512 453874 575572 453934
rect 575632 453874 575692 453934
rect 575752 453874 575812 453934
rect 575872 453874 575932 453934
rect 575992 453874 576052 453934
rect 576112 453874 576172 453934
rect 576232 453874 576292 453934
rect 576352 453874 576412 453934
rect 576472 453874 576532 453934
rect 576592 453874 576652 453934
rect 576712 453874 576772 453934
rect 576832 453874 576892 453934
rect 576952 453874 577012 453934
rect 577072 453874 577132 453934
rect 577192 453874 577252 453934
rect 577312 453874 577372 453934
rect 577432 453874 577492 453934
rect 577552 453874 577612 453934
rect 577672 453874 582788 453934
rect 567562 453859 582788 453874
rect 514788 453814 582788 453859
rect 514788 453799 572332 453814
rect 514788 453739 562222 453799
rect 562282 453739 562342 453799
rect 562402 453739 562462 453799
rect 562522 453739 562582 453799
rect 562642 453739 562702 453799
rect 562762 453739 562822 453799
rect 562882 453739 562942 453799
rect 563002 453739 563062 453799
rect 563122 453739 563182 453799
rect 563242 453739 563302 453799
rect 563362 453739 563422 453799
rect 563482 453739 563542 453799
rect 563602 453739 563662 453799
rect 563722 453739 563782 453799
rect 563842 453739 563902 453799
rect 563962 453739 564022 453799
rect 564082 453739 564142 453799
rect 564202 453739 564262 453799
rect 564322 453739 564382 453799
rect 564442 453739 564502 453799
rect 564562 453739 564622 453799
rect 564682 453739 564742 453799
rect 564802 453739 564862 453799
rect 564922 453739 564982 453799
rect 565042 453739 565102 453799
rect 565162 453739 565222 453799
rect 565282 453739 565342 453799
rect 565402 453739 565462 453799
rect 565522 453739 565582 453799
rect 565642 453739 565702 453799
rect 565762 453739 565822 453799
rect 565882 453739 565942 453799
rect 566002 453739 566062 453799
rect 566122 453739 566182 453799
rect 566242 453739 566302 453799
rect 566362 453739 566422 453799
rect 566482 453739 566542 453799
rect 566602 453739 566662 453799
rect 566722 453739 566782 453799
rect 566842 453739 566902 453799
rect 566962 453739 567022 453799
rect 567082 453739 567142 453799
rect 567202 453739 567262 453799
rect 567322 453739 567382 453799
rect 567442 453739 567502 453799
rect 567562 453754 572332 453799
rect 572392 453754 572452 453814
rect 572512 453754 572572 453814
rect 572632 453754 572692 453814
rect 572752 453754 572812 453814
rect 572872 453754 572932 453814
rect 572992 453754 573052 453814
rect 573112 453754 573172 453814
rect 573232 453754 573292 453814
rect 573352 453754 573412 453814
rect 573472 453754 573532 453814
rect 573592 453754 573652 453814
rect 573712 453754 573772 453814
rect 573832 453754 573892 453814
rect 573952 453754 574012 453814
rect 574072 453754 574132 453814
rect 574192 453754 574252 453814
rect 574312 453754 574372 453814
rect 574432 453754 574492 453814
rect 574552 453754 574612 453814
rect 574672 453754 574732 453814
rect 574792 453754 574852 453814
rect 574912 453754 574972 453814
rect 575032 453754 575092 453814
rect 575152 453754 575212 453814
rect 575272 453754 575332 453814
rect 575392 453754 575452 453814
rect 575512 453754 575572 453814
rect 575632 453754 575692 453814
rect 575752 453754 575812 453814
rect 575872 453754 575932 453814
rect 575992 453754 576052 453814
rect 576112 453754 576172 453814
rect 576232 453754 576292 453814
rect 576352 453754 576412 453814
rect 576472 453754 576532 453814
rect 576592 453754 576652 453814
rect 576712 453754 576772 453814
rect 576832 453754 576892 453814
rect 576952 453754 577012 453814
rect 577072 453754 577132 453814
rect 577192 453754 577252 453814
rect 577312 453754 577372 453814
rect 577432 453754 577492 453814
rect 577552 453754 577612 453814
rect 577672 453754 582788 453814
rect 567562 453739 582788 453754
rect 514788 449830 582788 453739
rect 583520 453264 584800 453376
rect 583520 452082 584800 452194
rect 583520 450900 584800 451012
rect 514788 449718 584800 449830
rect 514788 438756 582788 449718
rect 536882 426452 578882 426928
rect 536882 426216 572772 426452
rect 573008 426216 573244 426452
rect 573480 426216 573716 426452
rect 573952 426216 574188 426452
rect 574424 426216 574660 426452
rect 574896 426216 575132 426452
rect 575368 426216 575604 426452
rect 575840 426216 576076 426452
rect 576312 426216 576548 426452
rect 576784 426216 577020 426452
rect 577256 426216 578882 426452
rect 536882 425980 578882 426216
rect 536882 425744 572772 425980
rect 573008 425744 573244 425980
rect 573480 425744 573716 425980
rect 573952 425744 574188 425980
rect 574424 425744 574660 425980
rect 574896 425744 575132 425980
rect 575368 425744 575604 425980
rect 575840 425744 576076 425980
rect 576312 425744 576548 425980
rect 576784 425744 577020 425980
rect 577256 425744 578882 425980
rect 536882 425508 578882 425744
rect 536882 425272 572772 425508
rect 573008 425272 573244 425508
rect 573480 425272 573716 425508
rect 573952 425272 574188 425508
rect 574424 425272 574660 425508
rect 574896 425272 575132 425508
rect 575368 425272 575604 425508
rect 575840 425272 576076 425508
rect 576312 425272 576548 425508
rect 576784 425272 577020 425508
rect 577256 425272 578882 425508
rect -800 425086 480 425198
rect 536882 425036 578882 425272
rect 536882 424800 572772 425036
rect 573008 424800 573244 425036
rect 573480 424800 573716 425036
rect 573952 424800 574188 425036
rect 574424 424800 574660 425036
rect 574896 424800 575132 425036
rect 575368 424800 575604 425036
rect 575840 424800 576076 425036
rect 576312 424800 576548 425036
rect 576784 424800 577020 425036
rect 577256 424800 578882 425036
rect 536882 424564 578882 424800
rect 536882 424328 572772 424564
rect 573008 424328 573244 424564
rect 573480 424328 573716 424564
rect 573952 424328 574188 424564
rect 574424 424328 574660 424564
rect 574896 424328 575132 424564
rect 575368 424328 575604 424564
rect 575840 424328 576076 424564
rect 576312 424328 576548 424564
rect 576784 424328 577020 424564
rect 577256 424328 578882 424564
rect 536882 424092 578882 424328
rect -800 423904 480 424016
rect 536882 423856 572772 424092
rect 573008 423856 573244 424092
rect 573480 423856 573716 424092
rect 573952 423856 574188 424092
rect 574424 423856 574660 424092
rect 574896 423856 575132 424092
rect 575368 423856 575604 424092
rect 575840 423856 576076 424092
rect 576312 423856 576548 424092
rect 576784 423856 577020 424092
rect 577256 423856 578882 424092
rect 536882 423620 578882 423856
rect 536882 423384 572772 423620
rect 573008 423384 573244 423620
rect 573480 423384 573716 423620
rect 573952 423384 574188 423620
rect 574424 423384 574660 423620
rect 574896 423384 575132 423620
rect 575368 423384 575604 423620
rect 575840 423384 576076 423620
rect 576312 423384 576548 423620
rect 576784 423384 577020 423620
rect 577256 423384 578882 423620
rect 536882 423148 578882 423384
rect 536882 422912 572772 423148
rect 573008 422912 573244 423148
rect 573480 422912 573716 423148
rect 573952 422912 574188 423148
rect 574424 422912 574660 423148
rect 574896 422912 575132 423148
rect 575368 422912 575604 423148
rect 575840 422912 576076 423148
rect 576312 422912 576548 423148
rect 576784 422912 577020 423148
rect 577256 422912 578882 423148
rect -800 422722 480 422834
rect 536882 422676 578882 422912
rect 536882 422440 572772 422676
rect 573008 422440 573244 422676
rect 573480 422440 573716 422676
rect 573952 422440 574188 422676
rect 574424 422440 574660 422676
rect 574896 422440 575132 422676
rect 575368 422440 575604 422676
rect 575840 422440 576076 422676
rect 576312 422440 576548 422676
rect 576784 422440 577020 422676
rect 577256 422440 578882 422676
rect 536882 422204 578882 422440
rect 536882 421968 572772 422204
rect 573008 421968 573244 422204
rect 573480 421968 573716 422204
rect 573952 421968 574188 422204
rect 574424 421968 574660 422204
rect 574896 421968 575132 422204
rect 575368 421968 575604 422204
rect 575840 421968 576076 422204
rect 576312 421968 576548 422204
rect 576784 421968 577020 422204
rect 577256 421968 578882 422204
rect 536882 421732 578882 421968
rect -800 421540 480 421652
rect 536882 421496 572772 421732
rect 573008 421496 573244 421732
rect 573480 421496 573716 421732
rect 573952 421496 574188 421732
rect 574424 421496 574660 421732
rect 574896 421496 575132 421732
rect 575368 421496 575604 421732
rect 575840 421496 576076 421732
rect 576312 421496 576548 421732
rect 576784 421496 577020 421732
rect 577256 421496 578882 421732
rect 536882 421260 578882 421496
rect 536882 421024 572772 421260
rect 573008 421024 573244 421260
rect 573480 421024 573716 421260
rect 573952 421024 574188 421260
rect 574424 421024 574660 421260
rect 574896 421024 575132 421260
rect 575368 421024 575604 421260
rect 575840 421024 576076 421260
rect 576312 421024 576548 421260
rect 576784 421024 577020 421260
rect 577256 421024 578882 421260
rect 536882 420788 578882 421024
rect 536882 420552 572772 420788
rect 573008 420552 573244 420788
rect 573480 420552 573716 420788
rect 573952 420552 574188 420788
rect 574424 420552 574660 420788
rect 574896 420552 575132 420788
rect 575368 420552 575604 420788
rect 575840 420552 576076 420788
rect 576312 420552 576548 420788
rect 576784 420552 577020 420788
rect 577256 420552 578882 420788
rect -800 420358 480 420470
rect 536882 420272 578882 420552
rect -800 419176 480 419288
rect 583520 411206 584800 411318
rect 583520 410024 584800 410136
rect 583520 408842 584800 408954
rect 583520 407660 584800 407772
rect 583520 406478 584800 406590
rect 583520 405296 584800 405408
rect -800 381864 480 381976
rect -800 380682 480 380794
rect -800 379500 480 379612
rect -800 378318 480 378430
rect 477192 377866 483800 378072
rect 477060 377836 567660 377866
rect 477060 377600 477192 377836
rect 477428 377600 477664 377836
rect 477900 377600 478136 377836
rect 478372 377600 478608 377836
rect 478844 377600 479080 377836
rect 479316 377600 479552 377836
rect 479788 377600 480024 377836
rect 480260 377600 480496 377836
rect 480732 377600 480968 377836
rect 481204 377600 481440 377836
rect 481676 377600 481912 377836
rect 482148 377600 482384 377836
rect 482620 377600 482856 377836
rect 483092 377600 483328 377836
rect 483564 377600 567660 377836
rect 477060 377364 562624 377600
rect 562860 377364 563096 377600
rect 563332 377364 563568 377600
rect 563804 377364 564040 377600
rect 564276 377364 564512 377600
rect 564748 377364 564984 377600
rect 565220 377364 565456 377600
rect 565692 377364 565928 377600
rect 566164 377364 566400 377600
rect 566636 377364 566872 377600
rect 567108 377364 567660 377600
rect -800 377136 480 377248
rect 477060 377128 477192 377364
rect 477428 377128 477664 377364
rect 477900 377128 478136 377364
rect 478372 377128 478608 377364
rect 478844 377128 479080 377364
rect 479316 377128 479552 377364
rect 479788 377128 480024 377364
rect 480260 377128 480496 377364
rect 480732 377128 480968 377364
rect 481204 377128 481440 377364
rect 481676 377128 481912 377364
rect 482148 377128 482384 377364
rect 482620 377128 482856 377364
rect 483092 377128 483328 377364
rect 483564 377128 567660 377364
rect 477060 376892 562624 377128
rect 562860 376892 563096 377128
rect 563332 376892 563568 377128
rect 563804 376892 564040 377128
rect 564276 376892 564512 377128
rect 564748 376892 564984 377128
rect 565220 376892 565456 377128
rect 565692 376892 565928 377128
rect 566164 376892 566400 377128
rect 566636 376892 566872 377128
rect 567108 376892 567660 377128
rect 477060 376656 477192 376892
rect 477428 376656 477664 376892
rect 477900 376656 478136 376892
rect 478372 376656 478608 376892
rect 478844 376656 479080 376892
rect 479316 376656 479552 376892
rect 479788 376656 480024 376892
rect 480260 376656 480496 376892
rect 480732 376656 480968 376892
rect 481204 376656 481440 376892
rect 481676 376656 481912 376892
rect 482148 376656 482384 376892
rect 482620 376656 482856 376892
rect 483092 376656 483328 376892
rect 483564 376656 567660 376892
rect 477060 376420 562624 376656
rect 562860 376420 563096 376656
rect 563332 376420 563568 376656
rect 563804 376420 564040 376656
rect 564276 376420 564512 376656
rect 564748 376420 564984 376656
rect 565220 376420 565456 376656
rect 565692 376420 565928 376656
rect 566164 376420 566400 376656
rect 566636 376420 566872 376656
rect 567108 376420 567660 376656
rect 477060 376184 477192 376420
rect 477428 376184 477664 376420
rect 477900 376184 478136 376420
rect 478372 376184 478608 376420
rect 478844 376184 479080 376420
rect 479316 376184 479552 376420
rect 479788 376184 480024 376420
rect 480260 376184 480496 376420
rect 480732 376184 480968 376420
rect 481204 376184 481440 376420
rect 481676 376184 481912 376420
rect 482148 376184 482384 376420
rect 482620 376184 482856 376420
rect 483092 376184 483328 376420
rect 483564 376184 567660 376420
rect -800 375954 480 376066
rect 477060 375948 562624 376184
rect 562860 375948 563096 376184
rect 563332 375948 563568 376184
rect 563804 375948 564040 376184
rect 564276 375948 564512 376184
rect 564748 375948 564984 376184
rect 565220 375948 565456 376184
rect 565692 375948 565928 376184
rect 566164 375948 566400 376184
rect 566636 375948 566872 376184
rect 567108 375948 567660 376184
rect 477060 375712 477192 375948
rect 477428 375712 477664 375948
rect 477900 375712 478136 375948
rect 478372 375712 478608 375948
rect 478844 375712 479080 375948
rect 479316 375712 479552 375948
rect 479788 375712 480024 375948
rect 480260 375712 480496 375948
rect 480732 375712 480968 375948
rect 481204 375712 481440 375948
rect 481676 375712 481912 375948
rect 482148 375712 482384 375948
rect 482620 375712 482856 375948
rect 483092 375712 483328 375948
rect 483564 375712 567660 375948
rect 477060 375476 562624 375712
rect 562860 375476 563096 375712
rect 563332 375476 563568 375712
rect 563804 375476 564040 375712
rect 564276 375476 564512 375712
rect 564748 375476 564984 375712
rect 565220 375476 565456 375712
rect 565692 375476 565928 375712
rect 566164 375476 566400 375712
rect 566636 375476 566872 375712
rect 567108 375476 567660 375712
rect 477060 375240 477192 375476
rect 477428 375240 477664 375476
rect 477900 375240 478136 375476
rect 478372 375240 478608 375476
rect 478844 375240 479080 375476
rect 479316 375240 479552 375476
rect 479788 375240 480024 375476
rect 480260 375240 480496 375476
rect 480732 375240 480968 375476
rect 481204 375240 481440 375476
rect 481676 375240 481912 375476
rect 482148 375240 482384 375476
rect 482620 375240 482856 375476
rect 483092 375240 483328 375476
rect 483564 375240 567660 375476
rect 477060 375004 562624 375240
rect 562860 375004 563096 375240
rect 563332 375004 563568 375240
rect 563804 375004 564040 375240
rect 564276 375004 564512 375240
rect 564748 375004 564984 375240
rect 565220 375004 565456 375240
rect 565692 375004 565928 375240
rect 566164 375004 566400 375240
rect 566636 375004 566872 375240
rect 567108 375004 567660 375240
rect 477060 374768 477192 375004
rect 477428 374768 477664 375004
rect 477900 374768 478136 375004
rect 478372 374768 478608 375004
rect 478844 374768 479080 375004
rect 479316 374768 479552 375004
rect 479788 374768 480024 375004
rect 480260 374768 480496 375004
rect 480732 374768 480968 375004
rect 481204 374768 481440 375004
rect 481676 374768 481912 375004
rect 482148 374768 482384 375004
rect 482620 374768 482856 375004
rect 483092 374768 483328 375004
rect 483564 374768 567660 375004
rect 477060 374532 562624 374768
rect 562860 374532 563096 374768
rect 563332 374532 563568 374768
rect 563804 374532 564040 374768
rect 564276 374532 564512 374768
rect 564748 374532 564984 374768
rect 565220 374532 565456 374768
rect 565692 374532 565928 374768
rect 566164 374532 566400 374768
rect 566636 374532 566872 374768
rect 567108 374532 567660 374768
rect 477060 374296 477192 374532
rect 477428 374296 477664 374532
rect 477900 374296 478136 374532
rect 478372 374296 478608 374532
rect 478844 374296 479080 374532
rect 479316 374296 479552 374532
rect 479788 374296 480024 374532
rect 480260 374296 480496 374532
rect 480732 374296 480968 374532
rect 481204 374296 481440 374532
rect 481676 374296 481912 374532
rect 482148 374296 482384 374532
rect 482620 374296 482856 374532
rect 483092 374296 483328 374532
rect 483564 374296 567660 374532
rect 477060 374060 562624 374296
rect 562860 374060 563096 374296
rect 563332 374060 563568 374296
rect 563804 374060 564040 374296
rect 564276 374060 564512 374296
rect 564748 374060 564984 374296
rect 565220 374060 565456 374296
rect 565692 374060 565928 374296
rect 566164 374060 566400 374296
rect 566636 374060 566872 374296
rect 567108 374060 567660 374296
rect 477060 373824 477192 374060
rect 477428 373824 477664 374060
rect 477900 373824 478136 374060
rect 478372 373824 478608 374060
rect 478844 373824 479080 374060
rect 479316 373824 479552 374060
rect 479788 373824 480024 374060
rect 480260 373824 480496 374060
rect 480732 373824 480968 374060
rect 481204 373824 481440 374060
rect 481676 373824 481912 374060
rect 482148 373824 482384 374060
rect 482620 373824 482856 374060
rect 483092 373824 483328 374060
rect 483564 373824 567660 374060
rect 477060 373588 562624 373824
rect 562860 373588 563096 373824
rect 563332 373588 563568 373824
rect 563804 373588 564040 373824
rect 564276 373588 564512 373824
rect 564748 373588 564984 373824
rect 565220 373588 565456 373824
rect 565692 373588 565928 373824
rect 566164 373588 566400 373824
rect 566636 373588 566872 373824
rect 567108 373588 567660 373824
rect 477060 373352 477192 373588
rect 477428 373352 477664 373588
rect 477900 373352 478136 373588
rect 478372 373352 478608 373588
rect 478844 373352 479080 373588
rect 479316 373352 479552 373588
rect 479788 373352 480024 373588
rect 480260 373352 480496 373588
rect 480732 373352 480968 373588
rect 481204 373352 481440 373588
rect 481676 373352 481912 373588
rect 482148 373352 482384 373588
rect 482620 373352 482856 373588
rect 483092 373352 483328 373588
rect 483564 373352 567660 373588
rect 477060 373116 562624 373352
rect 562860 373116 563096 373352
rect 563332 373116 563568 373352
rect 563804 373116 564040 373352
rect 564276 373116 564512 373352
rect 564748 373116 564984 373352
rect 565220 373116 565456 373352
rect 565692 373116 565928 373352
rect 566164 373116 566400 373352
rect 566636 373116 566872 373352
rect 567108 373116 567660 373352
rect 477060 372880 477192 373116
rect 477428 372880 477664 373116
rect 477900 372880 478136 373116
rect 478372 372880 478608 373116
rect 478844 372880 479080 373116
rect 479316 372880 479552 373116
rect 479788 372880 480024 373116
rect 480260 372880 480496 373116
rect 480732 372880 480968 373116
rect 481204 372880 481440 373116
rect 481676 372880 481912 373116
rect 482148 372880 482384 373116
rect 482620 372880 482856 373116
rect 483092 372880 483328 373116
rect 483564 372880 567660 373116
rect 477060 372644 562624 372880
rect 562860 372644 563096 372880
rect 563332 372644 563568 372880
rect 563804 372644 564040 372880
rect 564276 372644 564512 372880
rect 564748 372644 564984 372880
rect 565220 372644 565456 372880
rect 565692 372644 565928 372880
rect 566164 372644 566400 372880
rect 566636 372644 566872 372880
rect 567108 372644 567660 372880
rect 477060 372408 477192 372644
rect 477428 372408 477664 372644
rect 477900 372408 478136 372644
rect 478372 372408 478608 372644
rect 478844 372408 479080 372644
rect 479316 372408 479552 372644
rect 479788 372408 480024 372644
rect 480260 372408 480496 372644
rect 480732 372408 480968 372644
rect 481204 372408 481440 372644
rect 481676 372408 481912 372644
rect 482148 372408 482384 372644
rect 482620 372408 482856 372644
rect 483092 372408 483328 372644
rect 483564 372408 567660 372644
rect 477060 372172 562624 372408
rect 562860 372172 563096 372408
rect 563332 372172 563568 372408
rect 563804 372172 564040 372408
rect 564276 372172 564512 372408
rect 564748 372172 564984 372408
rect 565220 372172 565456 372408
rect 565692 372172 565928 372408
rect 566164 372172 566400 372408
rect 566636 372172 566872 372408
rect 567108 372172 567660 372408
rect 477060 371936 477192 372172
rect 477428 371936 477664 372172
rect 477900 371936 478136 372172
rect 478372 371936 478608 372172
rect 478844 371936 479080 372172
rect 479316 371936 479552 372172
rect 479788 371936 480024 372172
rect 480260 371936 480496 372172
rect 480732 371936 480968 372172
rect 481204 371936 481440 372172
rect 481676 371936 481912 372172
rect 482148 371936 482384 372172
rect 482620 371936 482856 372172
rect 483092 371936 483328 372172
rect 483564 371936 567660 372172
rect 477060 371700 562624 371936
rect 562860 371700 563096 371936
rect 563332 371700 563568 371936
rect 563804 371700 564040 371936
rect 564276 371700 564512 371936
rect 564748 371700 564984 371936
rect 565220 371700 565456 371936
rect 565692 371700 565928 371936
rect 566164 371700 566400 371936
rect 566636 371700 566872 371936
rect 567108 371700 567660 371936
rect 477060 371464 477192 371700
rect 477428 371464 477664 371700
rect 477900 371464 478136 371700
rect 478372 371464 478608 371700
rect 478844 371464 479080 371700
rect 479316 371464 479552 371700
rect 479788 371464 480024 371700
rect 480260 371464 480496 371700
rect 480732 371464 480968 371700
rect 481204 371464 481440 371700
rect 481676 371464 481912 371700
rect 482148 371464 482384 371700
rect 482620 371464 482856 371700
rect 483092 371464 483328 371700
rect 483564 371464 567660 371700
rect 477060 371228 562624 371464
rect 562860 371228 563096 371464
rect 563332 371228 563568 371464
rect 563804 371228 564040 371464
rect 564276 371228 564512 371464
rect 564748 371228 564984 371464
rect 565220 371228 565456 371464
rect 565692 371228 565928 371464
rect 566164 371228 566400 371464
rect 566636 371228 566872 371464
rect 567108 371228 567660 371464
rect 477060 371200 567660 371228
rect 583520 364784 584800 364896
rect 583520 363602 584800 363714
rect 583520 362420 584800 362532
rect 583520 361238 584800 361350
rect 583520 360056 584800 360168
rect 583520 358874 584800 358986
rect -800 338642 480 338754
rect -800 337460 480 337572
rect -800 336278 480 336390
rect -800 335096 480 335208
rect -800 333914 480 334026
rect -800 332732 480 332844
rect 583520 319562 584800 319674
rect 583520 318380 584800 318492
rect 583520 317198 584800 317310
rect 583520 316016 584800 316128
rect 583520 314834 584800 314946
rect 583520 313652 584800 313764
rect -800 295420 480 295532
rect -800 294238 480 294350
rect -800 293056 480 293168
rect -800 291874 480 291986
rect -800 290692 480 290804
rect -800 289510 480 289622
rect 583520 275140 584800 275252
rect 583520 273958 584800 274070
rect 583520 272776 584800 272888
rect 583520 271594 584800 271706
rect 583520 270412 584800 270524
rect 583520 269230 584800 269342
rect -800 252398 480 252510
rect -800 251216 480 251328
rect -800 250034 480 250146
rect -800 248852 480 248964
rect -800 247670 480 247782
rect -800 246488 480 246600
rect 582340 235230 584800 240030
rect 582340 225230 584800 230030
rect -800 214888 1660 219688
rect -800 204888 1660 209688
rect 582340 191430 584800 196230
rect 582340 181430 584800 186230
rect -800 172888 1660 177688
rect -800 162888 1660 167688
rect 582340 146830 584800 151630
rect 582340 136830 584800 141630
rect -800 124776 480 124888
rect -800 123594 480 123706
rect -800 122412 480 122524
rect -800 121230 480 121342
rect -800 120048 480 120160
rect -800 118866 480 118978
rect 583520 95118 584800 95230
rect 583520 93936 584800 94048
rect 583520 92754 584800 92866
rect 583520 91572 584800 91684
rect -800 81554 480 81666
rect -800 80372 480 80484
rect -800 79190 480 79302
rect -800 78008 480 78120
rect -800 76826 480 76938
rect -800 75644 480 75756
rect 583520 50460 584800 50572
rect 583520 49278 584800 49390
rect 583520 48096 584800 48208
rect 583520 46914 584800 47026
rect -800 38332 480 38444
rect -800 37150 480 37262
rect -800 35968 480 36080
rect -800 34786 480 34898
rect -800 33604 480 33716
rect -800 32422 480 32534
rect 583520 24002 584800 24114
rect 583520 22820 584800 22932
rect 583520 21638 584800 21750
rect 583520 20456 584800 20568
rect 583520 19274 584800 19386
rect 583520 18092 584800 18204
rect -800 16910 480 17022
rect 583520 16910 584800 17022
rect -800 15728 480 15840
rect 583520 15728 584800 15840
rect -800 14546 480 14658
rect 583520 14546 584800 14658
rect -800 13364 480 13476
rect 583520 13364 584800 13476
rect -800 12182 480 12294
rect 583520 12182 584800 12294
rect -800 11000 480 11112
rect 583520 11000 584800 11112
rect -800 9818 480 9930
rect 583520 9818 584800 9930
rect -800 8636 480 8748
rect 583520 8636 584800 8748
rect -800 7454 480 7566
rect 583520 7454 584800 7566
rect -800 6272 480 6384
rect 583520 6272 584800 6384
rect -800 5090 480 5202
rect 583520 5090 584800 5202
rect -800 3908 480 4020
rect 583520 3908 584800 4020
rect -800 2726 480 2838
rect 583520 2726 584800 2838
rect -800 1544 480 1656
rect 583520 1544 584800 1656
<< via3 >>
rect 171000 692600 173000 697200
rect 173400 692600 175400 697200
rect 222706 692600 224706 697200
rect 225106 692600 227106 697200
rect 324412 692600 326412 697200
rect 326812 692600 328812 697200
rect 510654 692560 515334 697360
rect 520654 692560 525334 697360
rect 562600 639844 567400 644524
rect 562600 629844 567400 634524
rect 477192 522626 477428 522862
rect 477664 522626 477900 522862
rect 478136 522626 478372 522862
rect 478608 522626 478844 522862
rect 479080 522626 479316 522862
rect 479552 522626 479788 522862
rect 480024 522626 480260 522862
rect 480496 522626 480732 522862
rect 480968 522626 481204 522862
rect 481440 522626 481676 522862
rect 481912 522626 482148 522862
rect 482384 522626 482620 522862
rect 482856 522626 483092 522862
rect 483328 522626 483564 522862
rect 562624 522504 562860 522740
rect 563096 522504 563332 522740
rect 563568 522504 563804 522740
rect 564040 522504 564276 522740
rect 564512 522504 564748 522740
rect 564984 522504 565220 522740
rect 565456 522504 565692 522740
rect 565928 522504 566164 522740
rect 566400 522504 566636 522740
rect 566872 522504 567108 522740
rect 477192 522154 477428 522390
rect 477664 522154 477900 522390
rect 478136 522154 478372 522390
rect 478608 522154 478844 522390
rect 479080 522154 479316 522390
rect 479552 522154 479788 522390
rect 480024 522154 480260 522390
rect 480496 522154 480732 522390
rect 480968 522154 481204 522390
rect 481440 522154 481676 522390
rect 481912 522154 482148 522390
rect 482384 522154 482620 522390
rect 482856 522154 483092 522390
rect 483328 522154 483564 522390
rect 562624 522032 562860 522268
rect 563096 522032 563332 522268
rect 563568 522032 563804 522268
rect 564040 522032 564276 522268
rect 564512 522032 564748 522268
rect 564984 522032 565220 522268
rect 565456 522032 565692 522268
rect 565928 522032 566164 522268
rect 566400 522032 566636 522268
rect 566872 522032 567108 522268
rect 477192 521682 477428 521918
rect 477664 521682 477900 521918
rect 478136 521682 478372 521918
rect 478608 521682 478844 521918
rect 479080 521682 479316 521918
rect 479552 521682 479788 521918
rect 480024 521682 480260 521918
rect 480496 521682 480732 521918
rect 480968 521682 481204 521918
rect 481440 521682 481676 521918
rect 481912 521682 482148 521918
rect 482384 521682 482620 521918
rect 482856 521682 483092 521918
rect 483328 521682 483564 521918
rect 562624 521560 562860 521796
rect 563096 521560 563332 521796
rect 563568 521560 563804 521796
rect 564040 521560 564276 521796
rect 564512 521560 564748 521796
rect 564984 521560 565220 521796
rect 565456 521560 565692 521796
rect 565928 521560 566164 521796
rect 566400 521560 566636 521796
rect 566872 521560 567108 521796
rect 477192 521210 477428 521446
rect 477664 521210 477900 521446
rect 478136 521210 478372 521446
rect 478608 521210 478844 521446
rect 479080 521210 479316 521446
rect 479552 521210 479788 521446
rect 480024 521210 480260 521446
rect 480496 521210 480732 521446
rect 480968 521210 481204 521446
rect 481440 521210 481676 521446
rect 481912 521210 482148 521446
rect 482384 521210 482620 521446
rect 482856 521210 483092 521446
rect 483328 521210 483564 521446
rect 562624 521088 562860 521324
rect 563096 521088 563332 521324
rect 563568 521088 563804 521324
rect 564040 521088 564276 521324
rect 564512 521088 564748 521324
rect 564984 521088 565220 521324
rect 565456 521088 565692 521324
rect 565928 521088 566164 521324
rect 566400 521088 566636 521324
rect 566872 521088 567108 521324
rect 477192 520738 477428 520974
rect 477664 520738 477900 520974
rect 478136 520738 478372 520974
rect 478608 520738 478844 520974
rect 479080 520738 479316 520974
rect 479552 520738 479788 520974
rect 480024 520738 480260 520974
rect 480496 520738 480732 520974
rect 480968 520738 481204 520974
rect 481440 520738 481676 520974
rect 481912 520738 482148 520974
rect 482384 520738 482620 520974
rect 482856 520738 483092 520974
rect 483328 520738 483564 520974
rect 562624 520616 562860 520852
rect 563096 520616 563332 520852
rect 563568 520616 563804 520852
rect 564040 520616 564276 520852
rect 564512 520616 564748 520852
rect 564984 520616 565220 520852
rect 565456 520616 565692 520852
rect 565928 520616 566164 520852
rect 566400 520616 566636 520852
rect 566872 520616 567108 520852
rect 477192 520266 477428 520502
rect 477664 520266 477900 520502
rect 478136 520266 478372 520502
rect 478608 520266 478844 520502
rect 479080 520266 479316 520502
rect 479552 520266 479788 520502
rect 480024 520266 480260 520502
rect 480496 520266 480732 520502
rect 480968 520266 481204 520502
rect 481440 520266 481676 520502
rect 481912 520266 482148 520502
rect 482384 520266 482620 520502
rect 482856 520266 483092 520502
rect 483328 520266 483564 520502
rect 562624 520144 562860 520380
rect 563096 520144 563332 520380
rect 563568 520144 563804 520380
rect 564040 520144 564276 520380
rect 564512 520144 564748 520380
rect 564984 520144 565220 520380
rect 565456 520144 565692 520380
rect 565928 520144 566164 520380
rect 566400 520144 566636 520380
rect 566872 520144 567108 520380
rect 477192 519794 477428 520030
rect 477664 519794 477900 520030
rect 478136 519794 478372 520030
rect 478608 519794 478844 520030
rect 479080 519794 479316 520030
rect 479552 519794 479788 520030
rect 480024 519794 480260 520030
rect 480496 519794 480732 520030
rect 480968 519794 481204 520030
rect 481440 519794 481676 520030
rect 481912 519794 482148 520030
rect 482384 519794 482620 520030
rect 482856 519794 483092 520030
rect 483328 519794 483564 520030
rect 562624 519672 562860 519908
rect 563096 519672 563332 519908
rect 563568 519672 563804 519908
rect 564040 519672 564276 519908
rect 564512 519672 564748 519908
rect 564984 519672 565220 519908
rect 565456 519672 565692 519908
rect 565928 519672 566164 519908
rect 566400 519672 566636 519908
rect 566872 519672 567108 519908
rect 477192 519322 477428 519558
rect 477664 519322 477900 519558
rect 478136 519322 478372 519558
rect 478608 519322 478844 519558
rect 479080 519322 479316 519558
rect 479552 519322 479788 519558
rect 480024 519322 480260 519558
rect 480496 519322 480732 519558
rect 480968 519322 481204 519558
rect 481440 519322 481676 519558
rect 481912 519322 482148 519558
rect 482384 519322 482620 519558
rect 482856 519322 483092 519558
rect 483328 519322 483564 519558
rect 562624 519200 562860 519436
rect 563096 519200 563332 519436
rect 563568 519200 563804 519436
rect 564040 519200 564276 519436
rect 564512 519200 564748 519436
rect 564984 519200 565220 519436
rect 565456 519200 565692 519436
rect 565928 519200 566164 519436
rect 566400 519200 566636 519436
rect 566872 519200 567108 519436
rect 477192 518850 477428 519086
rect 477664 518850 477900 519086
rect 478136 518850 478372 519086
rect 478608 518850 478844 519086
rect 479080 518850 479316 519086
rect 479552 518850 479788 519086
rect 480024 518850 480260 519086
rect 480496 518850 480732 519086
rect 480968 518850 481204 519086
rect 481440 518850 481676 519086
rect 481912 518850 482148 519086
rect 482384 518850 482620 519086
rect 482856 518850 483092 519086
rect 483328 518850 483564 519086
rect 562624 518728 562860 518964
rect 563096 518728 563332 518964
rect 563568 518728 563804 518964
rect 564040 518728 564276 518964
rect 564512 518728 564748 518964
rect 564984 518728 565220 518964
rect 565456 518728 565692 518964
rect 565928 518728 566164 518964
rect 566400 518728 566636 518964
rect 566872 518728 567108 518964
rect 477192 518378 477428 518614
rect 477664 518378 477900 518614
rect 478136 518378 478372 518614
rect 478608 518378 478844 518614
rect 479080 518378 479316 518614
rect 479552 518378 479788 518614
rect 480024 518378 480260 518614
rect 480496 518378 480732 518614
rect 480968 518378 481204 518614
rect 481440 518378 481676 518614
rect 481912 518378 482148 518614
rect 482384 518378 482620 518614
rect 482856 518378 483092 518614
rect 483328 518378 483564 518614
rect 562624 518256 562860 518492
rect 563096 518256 563332 518492
rect 563568 518256 563804 518492
rect 564040 518256 564276 518492
rect 564512 518256 564748 518492
rect 564984 518256 565220 518492
rect 565456 518256 565692 518492
rect 565928 518256 566164 518492
rect 566400 518256 566636 518492
rect 566872 518256 567108 518492
rect 477192 517906 477428 518142
rect 477664 517906 477900 518142
rect 478136 517906 478372 518142
rect 478608 517906 478844 518142
rect 479080 517906 479316 518142
rect 479552 517906 479788 518142
rect 480024 517906 480260 518142
rect 480496 517906 480732 518142
rect 480968 517906 481204 518142
rect 481440 517906 481676 518142
rect 481912 517906 482148 518142
rect 482384 517906 482620 518142
rect 482856 517906 483092 518142
rect 483328 517906 483564 518142
rect 562624 517784 562860 518020
rect 563096 517784 563332 518020
rect 563568 517784 563804 518020
rect 564040 517784 564276 518020
rect 564512 517784 564748 518020
rect 564984 517784 565220 518020
rect 565456 517784 565692 518020
rect 565928 517784 566164 518020
rect 566400 517784 566636 518020
rect 566872 517784 567108 518020
rect 477192 517434 477428 517670
rect 477664 517434 477900 517670
rect 478136 517434 478372 517670
rect 478608 517434 478844 517670
rect 479080 517434 479316 517670
rect 479552 517434 479788 517670
rect 480024 517434 480260 517670
rect 480496 517434 480732 517670
rect 480968 517434 481204 517670
rect 481440 517434 481676 517670
rect 481912 517434 482148 517670
rect 482384 517434 482620 517670
rect 482856 517434 483092 517670
rect 483328 517434 483564 517670
rect 562624 517312 562860 517548
rect 563096 517312 563332 517548
rect 563568 517312 563804 517548
rect 564040 517312 564276 517548
rect 564512 517312 564748 517548
rect 564984 517312 565220 517548
rect 565456 517312 565692 517548
rect 565928 517312 566164 517548
rect 566400 517312 566636 517548
rect 566872 517312 567108 517548
rect 477192 516962 477428 517198
rect 477664 516962 477900 517198
rect 478136 516962 478372 517198
rect 478608 516962 478844 517198
rect 479080 516962 479316 517198
rect 479552 516962 479788 517198
rect 480024 516962 480260 517198
rect 480496 516962 480732 517198
rect 480968 516962 481204 517198
rect 481440 516962 481676 517198
rect 481912 516962 482148 517198
rect 482384 516962 482620 517198
rect 482856 516962 483092 517198
rect 483328 516962 483564 517198
rect 562624 516840 562860 517076
rect 563096 516840 563332 517076
rect 563568 516840 563804 517076
rect 564040 516840 564276 517076
rect 564512 516840 564748 517076
rect 564984 516840 565220 517076
rect 565456 516840 565692 517076
rect 565928 516840 566164 517076
rect 566400 516840 566636 517076
rect 566872 516840 567108 517076
rect 477192 516490 477428 516726
rect 477664 516490 477900 516726
rect 478136 516490 478372 516726
rect 478608 516490 478844 516726
rect 479080 516490 479316 516726
rect 479552 516490 479788 516726
rect 480024 516490 480260 516726
rect 480496 516490 480732 516726
rect 480968 516490 481204 516726
rect 481440 516490 481676 516726
rect 481912 516490 482148 516726
rect 482384 516490 482620 516726
rect 482856 516490 483092 516726
rect 483328 516490 483564 516726
rect 562624 516368 562860 516604
rect 563096 516368 563332 516604
rect 563568 516368 563804 516604
rect 564040 516368 564276 516604
rect 564512 516368 564748 516604
rect 564984 516368 565220 516604
rect 565456 516368 565692 516604
rect 565928 516368 566164 516604
rect 566400 516368 566636 516604
rect 566872 516368 567108 516604
rect 562480 495662 562560 495742
rect 562640 495662 562720 495742
rect 562800 495662 562880 495742
rect 562960 495662 563040 495742
rect 563120 495662 563200 495742
rect 563280 495662 563360 495742
rect 563440 495662 563520 495742
rect 563600 495662 563680 495742
rect 563760 495662 563840 495742
rect 563920 495662 564000 495742
rect 564080 495662 564160 495742
rect 564240 495662 564320 495742
rect 564400 495662 564480 495742
rect 564560 495662 564640 495742
rect 564720 495662 564800 495742
rect 564880 495662 564960 495742
rect 565040 495662 565120 495742
rect 565200 495662 565280 495742
rect 565360 495662 565440 495742
rect 565520 495662 565600 495742
rect 565680 495662 565760 495742
rect 565840 495662 565920 495742
rect 566000 495662 566080 495742
rect 566160 495662 566240 495742
rect 566320 495662 566400 495742
rect 566480 495662 566560 495742
rect 566640 495662 566720 495742
rect 566800 495662 566880 495742
rect 566960 495662 567040 495742
rect 567120 495662 567200 495742
rect 567280 495662 567360 495742
rect 562480 495502 562560 495582
rect 562640 495502 562720 495582
rect 562800 495502 562880 495582
rect 562960 495502 563040 495582
rect 563120 495502 563200 495582
rect 563280 495502 563360 495582
rect 563440 495502 563520 495582
rect 563600 495502 563680 495582
rect 563760 495502 563840 495582
rect 563920 495502 564000 495582
rect 564080 495502 564160 495582
rect 564240 495502 564320 495582
rect 564400 495502 564480 495582
rect 564560 495502 564640 495582
rect 564720 495502 564800 495582
rect 564880 495502 564960 495582
rect 565040 495502 565120 495582
rect 565200 495502 565280 495582
rect 565360 495502 565440 495582
rect 565520 495502 565600 495582
rect 565680 495502 565760 495582
rect 565840 495502 565920 495582
rect 566000 495502 566080 495582
rect 566160 495502 566240 495582
rect 566320 495502 566400 495582
rect 566480 495502 566560 495582
rect 566640 495502 566720 495582
rect 566800 495502 566880 495582
rect 566960 495502 567040 495582
rect 567120 495502 567200 495582
rect 567280 495502 567360 495582
rect 572640 495662 572720 495742
rect 572800 495662 572880 495742
rect 572960 495662 573040 495742
rect 573120 495662 573200 495742
rect 573280 495662 573360 495742
rect 573440 495662 573520 495742
rect 573600 495662 573680 495742
rect 573760 495662 573840 495742
rect 573920 495662 574000 495742
rect 574080 495662 574160 495742
rect 574240 495662 574320 495742
rect 574400 495662 574480 495742
rect 574560 495662 574640 495742
rect 574720 495662 574800 495742
rect 574880 495662 574960 495742
rect 575040 495662 575120 495742
rect 575200 495662 575280 495742
rect 575360 495662 575440 495742
rect 575520 495662 575600 495742
rect 575680 495662 575760 495742
rect 575840 495662 575920 495742
rect 576000 495662 576080 495742
rect 576160 495662 576240 495742
rect 576320 495662 576400 495742
rect 576480 495662 576560 495742
rect 576640 495662 576720 495742
rect 576800 495662 576880 495742
rect 576960 495662 577040 495742
rect 577120 495662 577200 495742
rect 577280 495662 577360 495742
rect 577440 495662 577520 495742
rect 572640 495502 572720 495582
rect 572800 495502 572880 495582
rect 572960 495502 573040 495582
rect 573120 495502 573200 495582
rect 573280 495502 573360 495582
rect 573440 495502 573520 495582
rect 573600 495502 573680 495582
rect 573760 495502 573840 495582
rect 573920 495502 574000 495582
rect 574080 495502 574160 495582
rect 574240 495502 574320 495582
rect 574400 495502 574480 495582
rect 574560 495502 574640 495582
rect 574720 495502 574800 495582
rect 574880 495502 574960 495582
rect 575040 495502 575120 495582
rect 575200 495502 575280 495582
rect 575360 495502 575440 495582
rect 575520 495502 575600 495582
rect 575680 495502 575760 495582
rect 575840 495502 575920 495582
rect 576000 495502 576080 495582
rect 576160 495502 576240 495582
rect 576320 495502 576400 495582
rect 576480 495502 576560 495582
rect 576640 495502 576720 495582
rect 576800 495502 576880 495582
rect 576960 495502 577040 495582
rect 577120 495502 577200 495582
rect 577280 495502 577360 495582
rect 577440 495502 577520 495582
rect 511616 494464 511680 494528
rect 511744 494464 511808 494528
rect 511872 494464 511936 494528
rect 512000 494464 512064 494528
rect 511616 494336 511680 494400
rect 511744 494336 511808 494400
rect 511872 494336 511936 494400
rect 512000 494336 512064 494400
rect 511616 494208 511680 494272
rect 511744 494208 511808 494272
rect 511872 494208 511936 494272
rect 512000 494208 512064 494272
rect 511616 494080 511680 494144
rect 511744 494080 511808 494144
rect 511872 494080 511936 494144
rect 512000 494080 512064 494144
rect 511616 493952 511680 494016
rect 511744 493952 511808 494016
rect 511872 493952 511936 494016
rect 512000 493952 512064 494016
rect 511616 493824 511680 493888
rect 511744 493824 511808 493888
rect 511872 493824 511936 493888
rect 512000 493824 512064 493888
rect 572772 483564 573008 483800
rect 573244 483564 573480 483800
rect 573716 483564 573952 483800
rect 574188 483564 574424 483800
rect 574660 483564 574896 483800
rect 575132 483564 575368 483800
rect 575604 483564 575840 483800
rect 576076 483564 576312 483800
rect 576548 483564 576784 483800
rect 577020 483564 577256 483800
rect 572772 483092 573008 483328
rect 573244 483092 573480 483328
rect 573716 483092 573952 483328
rect 574188 483092 574424 483328
rect 574660 483092 574896 483328
rect 575132 483092 575368 483328
rect 575604 483092 575840 483328
rect 576076 483092 576312 483328
rect 576548 483092 576784 483328
rect 577020 483092 577256 483328
rect 572772 482620 573008 482856
rect 573244 482620 573480 482856
rect 573716 482620 573952 482856
rect 574188 482620 574424 482856
rect 574660 482620 574896 482856
rect 575132 482620 575368 482856
rect 575604 482620 575840 482856
rect 576076 482620 576312 482856
rect 576548 482620 576784 482856
rect 577020 482620 577256 482856
rect 572772 482148 573008 482384
rect 573244 482148 573480 482384
rect 573716 482148 573952 482384
rect 574188 482148 574424 482384
rect 574660 482148 574896 482384
rect 575132 482148 575368 482384
rect 575604 482148 575840 482384
rect 576076 482148 576312 482384
rect 576548 482148 576784 482384
rect 577020 482148 577256 482384
rect 572772 481676 573008 481912
rect 573244 481676 573480 481912
rect 573716 481676 573952 481912
rect 574188 481676 574424 481912
rect 574660 481676 574896 481912
rect 575132 481676 575368 481912
rect 575604 481676 575840 481912
rect 576076 481676 576312 481912
rect 576548 481676 576784 481912
rect 577020 481676 577256 481912
rect 572772 481204 573008 481440
rect 573244 481204 573480 481440
rect 573716 481204 573952 481440
rect 574188 481204 574424 481440
rect 574660 481204 574896 481440
rect 575132 481204 575368 481440
rect 575604 481204 575840 481440
rect 576076 481204 576312 481440
rect 576548 481204 576784 481440
rect 577020 481204 577256 481440
rect 572772 480732 573008 480968
rect 573244 480732 573480 480968
rect 573716 480732 573952 480968
rect 574188 480732 574424 480968
rect 574660 480732 574896 480968
rect 575132 480732 575368 480968
rect 575604 480732 575840 480968
rect 576076 480732 576312 480968
rect 576548 480732 576784 480968
rect 577020 480732 577256 480968
rect 572772 480260 573008 480496
rect 573244 480260 573480 480496
rect 573716 480260 573952 480496
rect 574188 480260 574424 480496
rect 574660 480260 574896 480496
rect 575132 480260 575368 480496
rect 575604 480260 575840 480496
rect 576076 480260 576312 480496
rect 576548 480260 576784 480496
rect 577020 480260 577256 480496
rect 572772 479788 573008 480024
rect 573244 479788 573480 480024
rect 573716 479788 573952 480024
rect 574188 479788 574424 480024
rect 574660 479788 574896 480024
rect 575132 479788 575368 480024
rect 575604 479788 575840 480024
rect 576076 479788 576312 480024
rect 576548 479788 576784 480024
rect 577020 479788 577256 480024
rect 572772 479316 573008 479552
rect 573244 479316 573480 479552
rect 573716 479316 573952 479552
rect 574188 479316 574424 479552
rect 574660 479316 574896 479552
rect 575132 479316 575368 479552
rect 575604 479316 575840 479552
rect 576076 479316 576312 479552
rect 576548 479316 576784 479552
rect 577020 479316 577256 479552
rect 572772 478844 573008 479080
rect 573244 478844 573480 479080
rect 573716 478844 573952 479080
rect 574188 478844 574424 479080
rect 574660 478844 574896 479080
rect 575132 478844 575368 479080
rect 575604 478844 575840 479080
rect 576076 478844 576312 479080
rect 576548 478844 576784 479080
rect 577020 478844 577256 479080
rect 572772 478372 573008 478608
rect 573244 478372 573480 478608
rect 573716 478372 573952 478608
rect 574188 478372 574424 478608
rect 574660 478372 574896 478608
rect 575132 478372 575368 478608
rect 575604 478372 575840 478608
rect 576076 478372 576312 478608
rect 576548 478372 576784 478608
rect 577020 478372 577256 478608
rect 572772 477900 573008 478136
rect 573244 477900 573480 478136
rect 573716 477900 573952 478136
rect 574188 477900 574424 478136
rect 574660 477900 574896 478136
rect 575132 477900 575368 478136
rect 575604 477900 575840 478136
rect 576076 477900 576312 478136
rect 576548 477900 576784 478136
rect 577020 477900 577256 478136
rect 562480 455360 562560 455440
rect 562640 455360 562720 455440
rect 562800 455360 562880 455440
rect 562960 455360 563040 455440
rect 563120 455360 563200 455440
rect 563280 455360 563360 455440
rect 563440 455360 563520 455440
rect 563600 455360 563680 455440
rect 563760 455360 563840 455440
rect 563920 455360 564000 455440
rect 564080 455360 564160 455440
rect 564240 455360 564320 455440
rect 564400 455360 564480 455440
rect 564560 455360 564640 455440
rect 564720 455360 564800 455440
rect 564880 455360 564960 455440
rect 565040 455360 565120 455440
rect 565200 455360 565280 455440
rect 565360 455360 565440 455440
rect 565520 455360 565600 455440
rect 565680 455360 565760 455440
rect 565840 455360 565920 455440
rect 566000 455360 566080 455440
rect 566160 455360 566240 455440
rect 566320 455360 566400 455440
rect 566480 455360 566560 455440
rect 566640 455360 566720 455440
rect 566800 455360 566880 455440
rect 566960 455360 567040 455440
rect 567120 455360 567200 455440
rect 567280 455360 567360 455440
rect 562480 455200 562560 455280
rect 562640 455200 562720 455280
rect 562800 455200 562880 455280
rect 562960 455200 563040 455280
rect 563120 455200 563200 455280
rect 563280 455200 563360 455280
rect 563440 455200 563520 455280
rect 563600 455200 563680 455280
rect 563760 455200 563840 455280
rect 563920 455200 564000 455280
rect 564080 455200 564160 455280
rect 564240 455200 564320 455280
rect 564400 455200 564480 455280
rect 564560 455200 564640 455280
rect 564720 455200 564800 455280
rect 564880 455200 564960 455280
rect 565040 455200 565120 455280
rect 565200 455200 565280 455280
rect 565360 455200 565440 455280
rect 565520 455200 565600 455280
rect 565680 455200 565760 455280
rect 565840 455200 565920 455280
rect 566000 455200 566080 455280
rect 566160 455200 566240 455280
rect 566320 455200 566400 455280
rect 566480 455200 566560 455280
rect 566640 455200 566720 455280
rect 566800 455200 566880 455280
rect 566960 455200 567040 455280
rect 567120 455200 567200 455280
rect 567280 455200 567360 455280
rect 572640 455360 572720 455440
rect 572800 455360 572880 455440
rect 572960 455360 573040 455440
rect 573120 455360 573200 455440
rect 573280 455360 573360 455440
rect 573440 455360 573520 455440
rect 573600 455360 573680 455440
rect 573760 455360 573840 455440
rect 573920 455360 574000 455440
rect 574080 455360 574160 455440
rect 574240 455360 574320 455440
rect 574400 455360 574480 455440
rect 574560 455360 574640 455440
rect 574720 455360 574800 455440
rect 574880 455360 574960 455440
rect 575040 455360 575120 455440
rect 575200 455360 575280 455440
rect 575360 455360 575440 455440
rect 575520 455360 575600 455440
rect 575680 455360 575760 455440
rect 575840 455360 575920 455440
rect 576000 455360 576080 455440
rect 576160 455360 576240 455440
rect 576320 455360 576400 455440
rect 576480 455360 576560 455440
rect 576640 455360 576720 455440
rect 576800 455360 576880 455440
rect 576960 455360 577040 455440
rect 577120 455360 577200 455440
rect 577280 455360 577360 455440
rect 577440 455360 577520 455440
rect 572640 455200 572720 455280
rect 572800 455200 572880 455280
rect 572960 455200 573040 455280
rect 573120 455200 573200 455280
rect 573280 455200 573360 455280
rect 573440 455200 573520 455280
rect 573600 455200 573680 455280
rect 573760 455200 573840 455280
rect 573920 455200 574000 455280
rect 574080 455200 574160 455280
rect 574240 455200 574320 455280
rect 574400 455200 574480 455280
rect 574560 455200 574640 455280
rect 574720 455200 574800 455280
rect 574880 455200 574960 455280
rect 575040 455200 575120 455280
rect 575200 455200 575280 455280
rect 575360 455200 575440 455280
rect 575520 455200 575600 455280
rect 575680 455200 575760 455280
rect 575840 455200 575920 455280
rect 576000 455200 576080 455280
rect 576160 455200 576240 455280
rect 576320 455200 576400 455280
rect 576480 455200 576560 455280
rect 576640 455200 576720 455280
rect 576800 455200 576880 455280
rect 576960 455200 577040 455280
rect 577120 455200 577200 455280
rect 577280 455200 577360 455280
rect 577440 455200 577520 455280
rect 572772 426216 573008 426452
rect 573244 426216 573480 426452
rect 573716 426216 573952 426452
rect 574188 426216 574424 426452
rect 574660 426216 574896 426452
rect 575132 426216 575368 426452
rect 575604 426216 575840 426452
rect 576076 426216 576312 426452
rect 576548 426216 576784 426452
rect 577020 426216 577256 426452
rect 572772 425744 573008 425980
rect 573244 425744 573480 425980
rect 573716 425744 573952 425980
rect 574188 425744 574424 425980
rect 574660 425744 574896 425980
rect 575132 425744 575368 425980
rect 575604 425744 575840 425980
rect 576076 425744 576312 425980
rect 576548 425744 576784 425980
rect 577020 425744 577256 425980
rect 572772 425272 573008 425508
rect 573244 425272 573480 425508
rect 573716 425272 573952 425508
rect 574188 425272 574424 425508
rect 574660 425272 574896 425508
rect 575132 425272 575368 425508
rect 575604 425272 575840 425508
rect 576076 425272 576312 425508
rect 576548 425272 576784 425508
rect 577020 425272 577256 425508
rect 572772 424800 573008 425036
rect 573244 424800 573480 425036
rect 573716 424800 573952 425036
rect 574188 424800 574424 425036
rect 574660 424800 574896 425036
rect 575132 424800 575368 425036
rect 575604 424800 575840 425036
rect 576076 424800 576312 425036
rect 576548 424800 576784 425036
rect 577020 424800 577256 425036
rect 572772 424328 573008 424564
rect 573244 424328 573480 424564
rect 573716 424328 573952 424564
rect 574188 424328 574424 424564
rect 574660 424328 574896 424564
rect 575132 424328 575368 424564
rect 575604 424328 575840 424564
rect 576076 424328 576312 424564
rect 576548 424328 576784 424564
rect 577020 424328 577256 424564
rect 572772 423856 573008 424092
rect 573244 423856 573480 424092
rect 573716 423856 573952 424092
rect 574188 423856 574424 424092
rect 574660 423856 574896 424092
rect 575132 423856 575368 424092
rect 575604 423856 575840 424092
rect 576076 423856 576312 424092
rect 576548 423856 576784 424092
rect 577020 423856 577256 424092
rect 572772 423384 573008 423620
rect 573244 423384 573480 423620
rect 573716 423384 573952 423620
rect 574188 423384 574424 423620
rect 574660 423384 574896 423620
rect 575132 423384 575368 423620
rect 575604 423384 575840 423620
rect 576076 423384 576312 423620
rect 576548 423384 576784 423620
rect 577020 423384 577256 423620
rect 572772 422912 573008 423148
rect 573244 422912 573480 423148
rect 573716 422912 573952 423148
rect 574188 422912 574424 423148
rect 574660 422912 574896 423148
rect 575132 422912 575368 423148
rect 575604 422912 575840 423148
rect 576076 422912 576312 423148
rect 576548 422912 576784 423148
rect 577020 422912 577256 423148
rect 572772 422440 573008 422676
rect 573244 422440 573480 422676
rect 573716 422440 573952 422676
rect 574188 422440 574424 422676
rect 574660 422440 574896 422676
rect 575132 422440 575368 422676
rect 575604 422440 575840 422676
rect 576076 422440 576312 422676
rect 576548 422440 576784 422676
rect 577020 422440 577256 422676
rect 572772 421968 573008 422204
rect 573244 421968 573480 422204
rect 573716 421968 573952 422204
rect 574188 421968 574424 422204
rect 574660 421968 574896 422204
rect 575132 421968 575368 422204
rect 575604 421968 575840 422204
rect 576076 421968 576312 422204
rect 576548 421968 576784 422204
rect 577020 421968 577256 422204
rect 572772 421496 573008 421732
rect 573244 421496 573480 421732
rect 573716 421496 573952 421732
rect 574188 421496 574424 421732
rect 574660 421496 574896 421732
rect 575132 421496 575368 421732
rect 575604 421496 575840 421732
rect 576076 421496 576312 421732
rect 576548 421496 576784 421732
rect 577020 421496 577256 421732
rect 572772 421024 573008 421260
rect 573244 421024 573480 421260
rect 573716 421024 573952 421260
rect 574188 421024 574424 421260
rect 574660 421024 574896 421260
rect 575132 421024 575368 421260
rect 575604 421024 575840 421260
rect 576076 421024 576312 421260
rect 576548 421024 576784 421260
rect 577020 421024 577256 421260
rect 572772 420552 573008 420788
rect 573244 420552 573480 420788
rect 573716 420552 573952 420788
rect 574188 420552 574424 420788
rect 574660 420552 574896 420788
rect 575132 420552 575368 420788
rect 575604 420552 575840 420788
rect 576076 420552 576312 420788
rect 576548 420552 576784 420788
rect 577020 420552 577256 420788
rect 477192 377600 477428 377836
rect 477664 377600 477900 377836
rect 478136 377600 478372 377836
rect 478608 377600 478844 377836
rect 479080 377600 479316 377836
rect 479552 377600 479788 377836
rect 480024 377600 480260 377836
rect 480496 377600 480732 377836
rect 480968 377600 481204 377836
rect 481440 377600 481676 377836
rect 481912 377600 482148 377836
rect 482384 377600 482620 377836
rect 482856 377600 483092 377836
rect 483328 377600 483564 377836
rect 562624 377364 562860 377600
rect 563096 377364 563332 377600
rect 563568 377364 563804 377600
rect 564040 377364 564276 377600
rect 564512 377364 564748 377600
rect 564984 377364 565220 377600
rect 565456 377364 565692 377600
rect 565928 377364 566164 377600
rect 566400 377364 566636 377600
rect 566872 377364 567108 377600
rect 477192 377128 477428 377364
rect 477664 377128 477900 377364
rect 478136 377128 478372 377364
rect 478608 377128 478844 377364
rect 479080 377128 479316 377364
rect 479552 377128 479788 377364
rect 480024 377128 480260 377364
rect 480496 377128 480732 377364
rect 480968 377128 481204 377364
rect 481440 377128 481676 377364
rect 481912 377128 482148 377364
rect 482384 377128 482620 377364
rect 482856 377128 483092 377364
rect 483328 377128 483564 377364
rect 562624 376892 562860 377128
rect 563096 376892 563332 377128
rect 563568 376892 563804 377128
rect 564040 376892 564276 377128
rect 564512 376892 564748 377128
rect 564984 376892 565220 377128
rect 565456 376892 565692 377128
rect 565928 376892 566164 377128
rect 566400 376892 566636 377128
rect 566872 376892 567108 377128
rect 477192 376656 477428 376892
rect 477664 376656 477900 376892
rect 478136 376656 478372 376892
rect 478608 376656 478844 376892
rect 479080 376656 479316 376892
rect 479552 376656 479788 376892
rect 480024 376656 480260 376892
rect 480496 376656 480732 376892
rect 480968 376656 481204 376892
rect 481440 376656 481676 376892
rect 481912 376656 482148 376892
rect 482384 376656 482620 376892
rect 482856 376656 483092 376892
rect 483328 376656 483564 376892
rect 562624 376420 562860 376656
rect 563096 376420 563332 376656
rect 563568 376420 563804 376656
rect 564040 376420 564276 376656
rect 564512 376420 564748 376656
rect 564984 376420 565220 376656
rect 565456 376420 565692 376656
rect 565928 376420 566164 376656
rect 566400 376420 566636 376656
rect 566872 376420 567108 376656
rect 477192 376184 477428 376420
rect 477664 376184 477900 376420
rect 478136 376184 478372 376420
rect 478608 376184 478844 376420
rect 479080 376184 479316 376420
rect 479552 376184 479788 376420
rect 480024 376184 480260 376420
rect 480496 376184 480732 376420
rect 480968 376184 481204 376420
rect 481440 376184 481676 376420
rect 481912 376184 482148 376420
rect 482384 376184 482620 376420
rect 482856 376184 483092 376420
rect 483328 376184 483564 376420
rect 562624 375948 562860 376184
rect 563096 375948 563332 376184
rect 563568 375948 563804 376184
rect 564040 375948 564276 376184
rect 564512 375948 564748 376184
rect 564984 375948 565220 376184
rect 565456 375948 565692 376184
rect 565928 375948 566164 376184
rect 566400 375948 566636 376184
rect 566872 375948 567108 376184
rect 477192 375712 477428 375948
rect 477664 375712 477900 375948
rect 478136 375712 478372 375948
rect 478608 375712 478844 375948
rect 479080 375712 479316 375948
rect 479552 375712 479788 375948
rect 480024 375712 480260 375948
rect 480496 375712 480732 375948
rect 480968 375712 481204 375948
rect 481440 375712 481676 375948
rect 481912 375712 482148 375948
rect 482384 375712 482620 375948
rect 482856 375712 483092 375948
rect 483328 375712 483564 375948
rect 562624 375476 562860 375712
rect 563096 375476 563332 375712
rect 563568 375476 563804 375712
rect 564040 375476 564276 375712
rect 564512 375476 564748 375712
rect 564984 375476 565220 375712
rect 565456 375476 565692 375712
rect 565928 375476 566164 375712
rect 566400 375476 566636 375712
rect 566872 375476 567108 375712
rect 477192 375240 477428 375476
rect 477664 375240 477900 375476
rect 478136 375240 478372 375476
rect 478608 375240 478844 375476
rect 479080 375240 479316 375476
rect 479552 375240 479788 375476
rect 480024 375240 480260 375476
rect 480496 375240 480732 375476
rect 480968 375240 481204 375476
rect 481440 375240 481676 375476
rect 481912 375240 482148 375476
rect 482384 375240 482620 375476
rect 482856 375240 483092 375476
rect 483328 375240 483564 375476
rect 562624 375004 562860 375240
rect 563096 375004 563332 375240
rect 563568 375004 563804 375240
rect 564040 375004 564276 375240
rect 564512 375004 564748 375240
rect 564984 375004 565220 375240
rect 565456 375004 565692 375240
rect 565928 375004 566164 375240
rect 566400 375004 566636 375240
rect 566872 375004 567108 375240
rect 477192 374768 477428 375004
rect 477664 374768 477900 375004
rect 478136 374768 478372 375004
rect 478608 374768 478844 375004
rect 479080 374768 479316 375004
rect 479552 374768 479788 375004
rect 480024 374768 480260 375004
rect 480496 374768 480732 375004
rect 480968 374768 481204 375004
rect 481440 374768 481676 375004
rect 481912 374768 482148 375004
rect 482384 374768 482620 375004
rect 482856 374768 483092 375004
rect 483328 374768 483564 375004
rect 562624 374532 562860 374768
rect 563096 374532 563332 374768
rect 563568 374532 563804 374768
rect 564040 374532 564276 374768
rect 564512 374532 564748 374768
rect 564984 374532 565220 374768
rect 565456 374532 565692 374768
rect 565928 374532 566164 374768
rect 566400 374532 566636 374768
rect 566872 374532 567108 374768
rect 477192 374296 477428 374532
rect 477664 374296 477900 374532
rect 478136 374296 478372 374532
rect 478608 374296 478844 374532
rect 479080 374296 479316 374532
rect 479552 374296 479788 374532
rect 480024 374296 480260 374532
rect 480496 374296 480732 374532
rect 480968 374296 481204 374532
rect 481440 374296 481676 374532
rect 481912 374296 482148 374532
rect 482384 374296 482620 374532
rect 482856 374296 483092 374532
rect 483328 374296 483564 374532
rect 562624 374060 562860 374296
rect 563096 374060 563332 374296
rect 563568 374060 563804 374296
rect 564040 374060 564276 374296
rect 564512 374060 564748 374296
rect 564984 374060 565220 374296
rect 565456 374060 565692 374296
rect 565928 374060 566164 374296
rect 566400 374060 566636 374296
rect 566872 374060 567108 374296
rect 477192 373824 477428 374060
rect 477664 373824 477900 374060
rect 478136 373824 478372 374060
rect 478608 373824 478844 374060
rect 479080 373824 479316 374060
rect 479552 373824 479788 374060
rect 480024 373824 480260 374060
rect 480496 373824 480732 374060
rect 480968 373824 481204 374060
rect 481440 373824 481676 374060
rect 481912 373824 482148 374060
rect 482384 373824 482620 374060
rect 482856 373824 483092 374060
rect 483328 373824 483564 374060
rect 562624 373588 562860 373824
rect 563096 373588 563332 373824
rect 563568 373588 563804 373824
rect 564040 373588 564276 373824
rect 564512 373588 564748 373824
rect 564984 373588 565220 373824
rect 565456 373588 565692 373824
rect 565928 373588 566164 373824
rect 566400 373588 566636 373824
rect 566872 373588 567108 373824
rect 477192 373352 477428 373588
rect 477664 373352 477900 373588
rect 478136 373352 478372 373588
rect 478608 373352 478844 373588
rect 479080 373352 479316 373588
rect 479552 373352 479788 373588
rect 480024 373352 480260 373588
rect 480496 373352 480732 373588
rect 480968 373352 481204 373588
rect 481440 373352 481676 373588
rect 481912 373352 482148 373588
rect 482384 373352 482620 373588
rect 482856 373352 483092 373588
rect 483328 373352 483564 373588
rect 562624 373116 562860 373352
rect 563096 373116 563332 373352
rect 563568 373116 563804 373352
rect 564040 373116 564276 373352
rect 564512 373116 564748 373352
rect 564984 373116 565220 373352
rect 565456 373116 565692 373352
rect 565928 373116 566164 373352
rect 566400 373116 566636 373352
rect 566872 373116 567108 373352
rect 477192 372880 477428 373116
rect 477664 372880 477900 373116
rect 478136 372880 478372 373116
rect 478608 372880 478844 373116
rect 479080 372880 479316 373116
rect 479552 372880 479788 373116
rect 480024 372880 480260 373116
rect 480496 372880 480732 373116
rect 480968 372880 481204 373116
rect 481440 372880 481676 373116
rect 481912 372880 482148 373116
rect 482384 372880 482620 373116
rect 482856 372880 483092 373116
rect 483328 372880 483564 373116
rect 562624 372644 562860 372880
rect 563096 372644 563332 372880
rect 563568 372644 563804 372880
rect 564040 372644 564276 372880
rect 564512 372644 564748 372880
rect 564984 372644 565220 372880
rect 565456 372644 565692 372880
rect 565928 372644 566164 372880
rect 566400 372644 566636 372880
rect 566872 372644 567108 372880
rect 477192 372408 477428 372644
rect 477664 372408 477900 372644
rect 478136 372408 478372 372644
rect 478608 372408 478844 372644
rect 479080 372408 479316 372644
rect 479552 372408 479788 372644
rect 480024 372408 480260 372644
rect 480496 372408 480732 372644
rect 480968 372408 481204 372644
rect 481440 372408 481676 372644
rect 481912 372408 482148 372644
rect 482384 372408 482620 372644
rect 482856 372408 483092 372644
rect 483328 372408 483564 372644
rect 562624 372172 562860 372408
rect 563096 372172 563332 372408
rect 563568 372172 563804 372408
rect 564040 372172 564276 372408
rect 564512 372172 564748 372408
rect 564984 372172 565220 372408
rect 565456 372172 565692 372408
rect 565928 372172 566164 372408
rect 566400 372172 566636 372408
rect 566872 372172 567108 372408
rect 477192 371936 477428 372172
rect 477664 371936 477900 372172
rect 478136 371936 478372 372172
rect 478608 371936 478844 372172
rect 479080 371936 479316 372172
rect 479552 371936 479788 372172
rect 480024 371936 480260 372172
rect 480496 371936 480732 372172
rect 480968 371936 481204 372172
rect 481440 371936 481676 372172
rect 481912 371936 482148 372172
rect 482384 371936 482620 372172
rect 482856 371936 483092 372172
rect 483328 371936 483564 372172
rect 562624 371700 562860 371936
rect 563096 371700 563332 371936
rect 563568 371700 563804 371936
rect 564040 371700 564276 371936
rect 564512 371700 564748 371936
rect 564984 371700 565220 371936
rect 565456 371700 565692 371936
rect 565928 371700 566164 371936
rect 566400 371700 566636 371936
rect 566872 371700 567108 371936
rect 477192 371464 477428 371700
rect 477664 371464 477900 371700
rect 478136 371464 478372 371700
rect 478608 371464 478844 371700
rect 479080 371464 479316 371700
rect 479552 371464 479788 371700
rect 480024 371464 480260 371700
rect 480496 371464 480732 371700
rect 480968 371464 481204 371700
rect 481440 371464 481676 371700
rect 481912 371464 482148 371700
rect 482384 371464 482620 371700
rect 482856 371464 483092 371700
rect 483328 371464 483564 371700
rect 562624 371228 562860 371464
rect 563096 371228 563332 371464
rect 563568 371228 563804 371464
rect 564040 371228 564276 371464
rect 564512 371228 564748 371464
rect 564984 371228 565220 371464
rect 565456 371228 565692 371464
rect 565928 371228 566164 371464
rect 566400 371228 566636 371464
rect 566872 371228 567108 371464
<< metal4 >>
rect 115334 697380 577480 697420
rect 115334 697360 577492 697380
rect 115334 697200 510654 697360
rect 115334 692600 171000 697200
rect 173000 692600 173400 697200
rect 175400 692600 222706 697200
rect 224706 692600 225106 697200
rect 227106 692600 324412 697200
rect 326412 692600 326812 697200
rect 328812 692600 510654 697200
rect 115334 692560 510654 692600
rect 515334 692560 520654 697360
rect 525334 697144 577492 697360
rect 525334 696908 572772 697144
rect 573008 696908 573244 697144
rect 573480 696908 573716 697144
rect 573952 696908 574188 697144
rect 574424 696908 574660 697144
rect 574896 696908 575132 697144
rect 575368 696908 575604 697144
rect 575840 696908 576076 697144
rect 576312 696908 576548 697144
rect 576784 696908 577020 697144
rect 577256 696908 577492 697144
rect 525334 696672 577492 696908
rect 525334 696436 572772 696672
rect 573008 696436 573244 696672
rect 573480 696436 573716 696672
rect 573952 696436 574188 696672
rect 574424 696436 574660 696672
rect 574896 696436 575132 696672
rect 575368 696436 575604 696672
rect 575840 696436 576076 696672
rect 576312 696436 576548 696672
rect 576784 696436 577020 696672
rect 577256 696436 577492 696672
rect 525334 696200 577492 696436
rect 525334 695964 572772 696200
rect 573008 695964 573244 696200
rect 573480 695964 573716 696200
rect 573952 695964 574188 696200
rect 574424 695964 574660 696200
rect 574896 695964 575132 696200
rect 575368 695964 575604 696200
rect 575840 695964 576076 696200
rect 576312 695964 576548 696200
rect 576784 695964 577020 696200
rect 577256 695964 577492 696200
rect 525334 695728 577492 695964
rect 525334 695492 572772 695728
rect 573008 695492 573244 695728
rect 573480 695492 573716 695728
rect 573952 695492 574188 695728
rect 574424 695492 574660 695728
rect 574896 695492 575132 695728
rect 575368 695492 575604 695728
rect 575840 695492 576076 695728
rect 576312 695492 576548 695728
rect 576784 695492 577020 695728
rect 577256 695492 577492 695728
rect 525334 695256 577492 695492
rect 525334 695020 572772 695256
rect 573008 695020 573244 695256
rect 573480 695020 573716 695256
rect 573952 695020 574188 695256
rect 574424 695020 574660 695256
rect 574896 695020 575132 695256
rect 575368 695020 575604 695256
rect 575840 695020 576076 695256
rect 576312 695020 576548 695256
rect 576784 695020 577020 695256
rect 577256 695020 577492 695256
rect 525334 694784 577492 695020
rect 525334 694548 572772 694784
rect 573008 694548 573244 694784
rect 573480 694548 573716 694784
rect 573952 694548 574188 694784
rect 574424 694548 574660 694784
rect 574896 694548 575132 694784
rect 575368 694548 575604 694784
rect 575840 694548 576076 694784
rect 576312 694548 576548 694784
rect 576784 694548 577020 694784
rect 577256 694548 577492 694784
rect 525334 694312 577492 694548
rect 525334 694076 572772 694312
rect 573008 694076 573244 694312
rect 573480 694076 573716 694312
rect 573952 694076 574188 694312
rect 574424 694076 574660 694312
rect 574896 694076 575132 694312
rect 575368 694076 575604 694312
rect 575840 694076 576076 694312
rect 576312 694076 576548 694312
rect 576784 694076 577020 694312
rect 577256 694076 577492 694312
rect 525334 693840 577492 694076
rect 525334 693604 572772 693840
rect 573008 693604 573244 693840
rect 573480 693604 573716 693840
rect 573952 693604 574188 693840
rect 574424 693604 574660 693840
rect 574896 693604 575132 693840
rect 575368 693604 575604 693840
rect 575840 693604 576076 693840
rect 576312 693604 576548 693840
rect 576784 693604 577020 693840
rect 577256 693604 577492 693840
rect 525334 693368 577492 693604
rect 525334 693132 572772 693368
rect 573008 693132 573244 693368
rect 573480 693132 573716 693368
rect 573952 693132 574188 693368
rect 574424 693132 574660 693368
rect 574896 693132 575132 693368
rect 575368 693132 575604 693368
rect 575840 693132 576076 693368
rect 576312 693132 576548 693368
rect 576784 693132 577020 693368
rect 577256 693132 577492 693368
rect 525334 692896 577492 693132
rect 525334 692660 572772 692896
rect 573008 692660 573244 692896
rect 573480 692660 573716 692896
rect 573952 692660 574188 692896
rect 574424 692660 574660 692896
rect 574896 692660 575132 692896
rect 575368 692660 575604 692896
rect 575840 692660 576076 692896
rect 576312 692660 576548 692896
rect 576784 692660 577020 692896
rect 577256 692660 577492 692896
rect 525334 692560 577480 692660
rect 115334 692500 577480 692560
rect 562456 644584 567424 644608
rect 562456 639784 562480 644584
rect 567400 639784 567424 644584
rect 562456 639760 567424 639784
rect 562456 634584 567424 634608
rect 562456 629784 562480 634584
rect 567400 629784 567424 634584
rect 562456 629760 567424 629784
rect 572600 623400 577400 623588
rect 477192 522892 483800 523098
rect 477060 522862 483800 522892
rect 477060 522626 477192 522862
rect 477428 522626 477664 522862
rect 477900 522626 478136 522862
rect 478372 522626 478608 522862
rect 478844 522626 479080 522862
rect 479316 522626 479552 522862
rect 479788 522626 480024 522862
rect 480260 522626 480496 522862
rect 480732 522626 480968 522862
rect 481204 522626 481440 522862
rect 481676 522626 481912 522862
rect 482148 522626 482384 522862
rect 482620 522626 482856 522862
rect 483092 522626 483328 522862
rect 483564 522626 483800 522862
rect 477060 522390 483800 522626
rect 477060 522154 477192 522390
rect 477428 522154 477664 522390
rect 477900 522154 478136 522390
rect 478372 522154 478608 522390
rect 478844 522154 479080 522390
rect 479316 522154 479552 522390
rect 479788 522154 480024 522390
rect 480260 522154 480496 522390
rect 480732 522154 480968 522390
rect 481204 522154 481440 522390
rect 481676 522154 481912 522390
rect 482148 522154 482384 522390
rect 482620 522154 482856 522390
rect 483092 522154 483328 522390
rect 483564 522154 483800 522390
rect 477060 521918 483800 522154
rect 477060 521682 477192 521918
rect 477428 521682 477664 521918
rect 477900 521682 478136 521918
rect 478372 521682 478608 521918
rect 478844 521682 479080 521918
rect 479316 521682 479552 521918
rect 479788 521682 480024 521918
rect 480260 521682 480496 521918
rect 480732 521682 480968 521918
rect 481204 521682 481440 521918
rect 481676 521682 481912 521918
rect 482148 521682 482384 521918
rect 482620 521682 482856 521918
rect 483092 521682 483328 521918
rect 483564 521682 483800 521918
rect 477060 521446 483800 521682
rect 477060 521210 477192 521446
rect 477428 521210 477664 521446
rect 477900 521210 478136 521446
rect 478372 521210 478608 521446
rect 478844 521210 479080 521446
rect 479316 521210 479552 521446
rect 479788 521210 480024 521446
rect 480260 521210 480496 521446
rect 480732 521210 480968 521446
rect 481204 521210 481440 521446
rect 481676 521210 481912 521446
rect 482148 521210 482384 521446
rect 482620 521210 482856 521446
rect 483092 521210 483328 521446
rect 483564 521210 483800 521446
rect 477060 520974 483800 521210
rect 477060 520738 477192 520974
rect 477428 520738 477664 520974
rect 477900 520738 478136 520974
rect 478372 520738 478608 520974
rect 478844 520738 479080 520974
rect 479316 520738 479552 520974
rect 479788 520738 480024 520974
rect 480260 520738 480496 520974
rect 480732 520738 480968 520974
rect 481204 520738 481440 520974
rect 481676 520738 481912 520974
rect 482148 520738 482384 520974
rect 482620 520738 482856 520974
rect 483092 520738 483328 520974
rect 483564 520738 483800 520974
rect 477060 520502 483800 520738
rect 477060 520266 477192 520502
rect 477428 520266 477664 520502
rect 477900 520266 478136 520502
rect 478372 520266 478608 520502
rect 478844 520266 479080 520502
rect 479316 520266 479552 520502
rect 479788 520266 480024 520502
rect 480260 520266 480496 520502
rect 480732 520266 480968 520502
rect 481204 520266 481440 520502
rect 481676 520266 481912 520502
rect 482148 520266 482384 520502
rect 482620 520266 482856 520502
rect 483092 520266 483328 520502
rect 483564 520266 483800 520502
rect 477060 520030 483800 520266
rect 477060 519794 477192 520030
rect 477428 519794 477664 520030
rect 477900 519794 478136 520030
rect 478372 519794 478608 520030
rect 478844 519794 479080 520030
rect 479316 519794 479552 520030
rect 479788 519794 480024 520030
rect 480260 519794 480496 520030
rect 480732 519794 480968 520030
rect 481204 519794 481440 520030
rect 481676 519794 481912 520030
rect 482148 519794 482384 520030
rect 482620 519794 482856 520030
rect 483092 519794 483328 520030
rect 483564 519794 483800 520030
rect 477060 519558 483800 519794
rect 477060 519322 477192 519558
rect 477428 519322 477664 519558
rect 477900 519322 478136 519558
rect 478372 519322 478608 519558
rect 478844 519322 479080 519558
rect 479316 519322 479552 519558
rect 479788 519322 480024 519558
rect 480260 519322 480496 519558
rect 480732 519322 480968 519558
rect 481204 519322 481440 519558
rect 481676 519322 481912 519558
rect 482148 519322 482384 519558
rect 482620 519322 482856 519558
rect 483092 519322 483328 519558
rect 483564 519322 483800 519558
rect 477060 519086 483800 519322
rect 477060 518850 477192 519086
rect 477428 518850 477664 519086
rect 477900 518850 478136 519086
rect 478372 518850 478608 519086
rect 478844 518850 479080 519086
rect 479316 518850 479552 519086
rect 479788 518850 480024 519086
rect 480260 518850 480496 519086
rect 480732 518850 480968 519086
rect 481204 518850 481440 519086
rect 481676 518850 481912 519086
rect 482148 518850 482384 519086
rect 482620 518850 482856 519086
rect 483092 518850 483328 519086
rect 483564 518850 483800 519086
rect 477060 518614 483800 518850
rect 477060 518378 477192 518614
rect 477428 518378 477664 518614
rect 477900 518378 478136 518614
rect 478372 518378 478608 518614
rect 478844 518378 479080 518614
rect 479316 518378 479552 518614
rect 479788 518378 480024 518614
rect 480260 518378 480496 518614
rect 480732 518378 480968 518614
rect 481204 518378 481440 518614
rect 481676 518378 481912 518614
rect 482148 518378 482384 518614
rect 482620 518378 482856 518614
rect 483092 518378 483328 518614
rect 483564 518378 483800 518614
rect 477060 518142 483800 518378
rect 477060 517906 477192 518142
rect 477428 517906 477664 518142
rect 477900 517906 478136 518142
rect 478372 517906 478608 518142
rect 478844 517906 479080 518142
rect 479316 517906 479552 518142
rect 479788 517906 480024 518142
rect 480260 517906 480496 518142
rect 480732 517906 480968 518142
rect 481204 517906 481440 518142
rect 481676 517906 481912 518142
rect 482148 517906 482384 518142
rect 482620 517906 482856 518142
rect 483092 517906 483328 518142
rect 483564 517906 483800 518142
rect 477060 517670 483800 517906
rect 477060 517434 477192 517670
rect 477428 517434 477664 517670
rect 477900 517434 478136 517670
rect 478372 517434 478608 517670
rect 478844 517434 479080 517670
rect 479316 517434 479552 517670
rect 479788 517434 480024 517670
rect 480260 517434 480496 517670
rect 480732 517434 480968 517670
rect 481204 517434 481440 517670
rect 481676 517434 481912 517670
rect 482148 517434 482384 517670
rect 482620 517434 482856 517670
rect 483092 517434 483328 517670
rect 483564 517434 483800 517670
rect 477060 517198 483800 517434
rect 477060 516962 477192 517198
rect 477428 516962 477664 517198
rect 477900 516962 478136 517198
rect 478372 516962 478608 517198
rect 478844 516962 479080 517198
rect 479316 516962 479552 517198
rect 479788 516962 480024 517198
rect 480260 516962 480496 517198
rect 480732 516962 480968 517198
rect 481204 516962 481440 517198
rect 481676 516962 481912 517198
rect 482148 516962 482384 517198
rect 482620 516962 482856 517198
rect 483092 516962 483328 517198
rect 483564 516962 483800 517198
rect 477060 516726 483800 516962
rect 477060 516490 477192 516726
rect 477428 516490 477664 516726
rect 477900 516490 478136 516726
rect 478372 516490 478608 516726
rect 478844 516490 479080 516726
rect 479316 516490 479552 516726
rect 479788 516490 480024 516726
rect 480260 516490 480496 516726
rect 480732 516490 480968 516726
rect 481204 516490 481440 516726
rect 481676 516490 481912 516726
rect 482148 516490 482384 516726
rect 482620 516490 482856 516726
rect 483092 516490 483328 516726
rect 483564 516490 483800 516726
rect 562388 522740 567816 523212
rect 477060 378072 483726 516490
rect 562388 516368 562624 522740
rect 562860 516368 563096 522740
rect 563332 516368 563568 522740
rect 563804 516368 564040 522740
rect 564276 516368 564512 522740
rect 564748 516368 564984 522740
rect 565220 516368 565456 522740
rect 565692 516368 565928 522740
rect 566164 516368 566400 522740
rect 566636 516368 566872 522740
rect 567108 516368 567816 522740
rect 562388 516132 567816 516368
rect 562380 495782 567480 495822
rect 562380 495742 562624 495782
rect 562860 495742 563096 495782
rect 563332 495742 563568 495782
rect 563804 495742 564040 495782
rect 564276 495742 564512 495782
rect 564748 495742 564984 495782
rect 565220 495742 565456 495782
rect 565692 495742 565928 495782
rect 566164 495742 566400 495782
rect 566636 495742 566872 495782
rect 567108 495742 567480 495782
rect 562380 495662 562480 495742
rect 562560 495662 562624 495742
rect 562880 495662 562960 495742
rect 563040 495662 563096 495742
rect 563360 495662 563440 495742
rect 563520 495662 563568 495742
rect 563840 495662 563920 495742
rect 564000 495662 564040 495742
rect 564320 495662 564400 495742
rect 564480 495662 564512 495742
rect 564800 495662 564880 495742
rect 564960 495662 564984 495742
rect 565280 495662 565360 495742
rect 565440 495662 565456 495742
rect 565760 495662 565840 495742
rect 565920 495662 565928 495742
rect 566240 495662 566320 495742
rect 566636 495662 566640 495742
rect 566720 495662 566800 495742
rect 567108 495662 567120 495742
rect 567200 495662 567280 495742
rect 567360 495662 567480 495742
rect 562380 495582 562624 495662
rect 562860 495582 563096 495662
rect 563332 495582 563568 495662
rect 563804 495582 564040 495662
rect 564276 495582 564512 495662
rect 564748 495582 564984 495662
rect 565220 495582 565456 495662
rect 565692 495582 565928 495662
rect 566164 495582 566400 495662
rect 566636 495582 566872 495662
rect 567108 495582 567480 495662
rect 562380 495502 562480 495582
rect 562560 495546 562624 495582
rect 562560 495502 562640 495546
rect 562720 495502 562800 495546
rect 562880 495502 562960 495582
rect 563040 495546 563096 495582
rect 563040 495502 563120 495546
rect 563200 495502 563280 495546
rect 563360 495502 563440 495582
rect 563520 495546 563568 495582
rect 563520 495502 563600 495546
rect 563680 495502 563760 495546
rect 563840 495502 563920 495582
rect 564000 495546 564040 495582
rect 564000 495502 564080 495546
rect 564160 495502 564240 495546
rect 564320 495502 564400 495582
rect 564480 495546 564512 495582
rect 564480 495502 564560 495546
rect 564640 495502 564720 495546
rect 564800 495502 564880 495582
rect 564960 495546 564984 495582
rect 564960 495502 565040 495546
rect 565120 495502 565200 495546
rect 565280 495502 565360 495582
rect 565440 495546 565456 495582
rect 565440 495502 565520 495546
rect 565600 495502 565680 495546
rect 565760 495502 565840 495582
rect 565920 495546 565928 495582
rect 565920 495502 566000 495546
rect 566080 495502 566160 495546
rect 566240 495502 566320 495582
rect 566636 495546 566640 495582
rect 566400 495502 566480 495546
rect 566560 495502 566640 495546
rect 566720 495502 566800 495582
rect 567108 495546 567120 495582
rect 566880 495502 566960 495546
rect 567040 495502 567120 495546
rect 567200 495502 567280 495582
rect 567360 495502 567480 495582
rect 562380 495462 567480 495502
rect 572540 495782 577640 495822
rect 572540 495742 572784 495782
rect 573020 495742 573256 495782
rect 573492 495742 573728 495782
rect 573964 495742 574200 495782
rect 574436 495742 574672 495782
rect 574908 495742 575144 495782
rect 575380 495742 575616 495782
rect 575852 495742 576088 495782
rect 576324 495742 576560 495782
rect 576796 495742 577032 495782
rect 577268 495742 577640 495782
rect 572540 495662 572640 495742
rect 572720 495662 572784 495742
rect 573040 495662 573120 495742
rect 573200 495662 573256 495742
rect 573520 495662 573600 495742
rect 573680 495662 573728 495742
rect 574000 495662 574080 495742
rect 574160 495662 574200 495742
rect 574480 495662 574560 495742
rect 574640 495662 574672 495742
rect 574960 495662 575040 495742
rect 575120 495662 575144 495742
rect 575440 495662 575520 495742
rect 575600 495662 575616 495742
rect 575920 495662 576000 495742
rect 576080 495662 576088 495742
rect 576400 495662 576480 495742
rect 576796 495662 576800 495742
rect 576880 495662 576960 495742
rect 577268 495662 577280 495742
rect 577360 495662 577440 495742
rect 577520 495662 577640 495742
rect 572540 495582 572784 495662
rect 573020 495582 573256 495662
rect 573492 495582 573728 495662
rect 573964 495582 574200 495662
rect 574436 495582 574672 495662
rect 574908 495582 575144 495662
rect 575380 495582 575616 495662
rect 575852 495582 576088 495662
rect 576324 495582 576560 495662
rect 576796 495582 577032 495662
rect 577268 495582 577640 495662
rect 572540 495502 572640 495582
rect 572720 495546 572784 495582
rect 572720 495502 572800 495546
rect 572880 495502 572960 495546
rect 573040 495502 573120 495582
rect 573200 495546 573256 495582
rect 573200 495502 573280 495546
rect 573360 495502 573440 495546
rect 573520 495502 573600 495582
rect 573680 495546 573728 495582
rect 573680 495502 573760 495546
rect 573840 495502 573920 495546
rect 574000 495502 574080 495582
rect 574160 495546 574200 495582
rect 574160 495502 574240 495546
rect 574320 495502 574400 495546
rect 574480 495502 574560 495582
rect 574640 495546 574672 495582
rect 574640 495502 574720 495546
rect 574800 495502 574880 495546
rect 574960 495502 575040 495582
rect 575120 495546 575144 495582
rect 575120 495502 575200 495546
rect 575280 495502 575360 495546
rect 575440 495502 575520 495582
rect 575600 495546 575616 495582
rect 575600 495502 575680 495546
rect 575760 495502 575840 495546
rect 575920 495502 576000 495582
rect 576080 495546 576088 495582
rect 576080 495502 576160 495546
rect 576240 495502 576320 495546
rect 576400 495502 576480 495582
rect 576796 495546 576800 495582
rect 576560 495502 576640 495546
rect 576720 495502 576800 495546
rect 576880 495502 576960 495582
rect 577268 495546 577280 495582
rect 577040 495502 577120 495546
rect 577200 495502 577280 495546
rect 577360 495502 577440 495582
rect 577520 495502 577640 495582
rect 572540 495462 577640 495502
rect 511584 494528 512160 494700
rect 511584 494464 511616 494528
rect 511680 494464 511744 494528
rect 511808 494464 511872 494528
rect 511936 494464 512000 494528
rect 512064 494464 512160 494528
rect 511584 494400 512160 494464
rect 511584 494336 511616 494400
rect 511680 494336 511744 494400
rect 511808 494336 511872 494400
rect 511936 494336 512000 494400
rect 512064 494336 512160 494400
rect 511584 494272 512160 494336
rect 511584 494208 511616 494272
rect 511680 494208 511744 494272
rect 511808 494208 511872 494272
rect 511936 494208 512000 494272
rect 512064 494208 512160 494272
rect 511584 494144 512160 494208
rect 511584 494080 511616 494144
rect 511680 494080 511744 494144
rect 511808 494080 511872 494144
rect 511936 494080 512000 494144
rect 512064 494080 512160 494144
rect 511584 494016 512160 494080
rect 511584 493952 511616 494016
rect 511680 493952 511744 494016
rect 511808 493952 511872 494016
rect 511936 493952 512000 494016
rect 512064 493952 512160 494016
rect 511584 493888 512160 493952
rect 511584 493824 511616 493888
rect 511680 493824 511744 493888
rect 511808 493824 511872 493888
rect 511936 493824 512000 493888
rect 512064 493824 512160 493888
rect 511584 475300 512160 493824
rect 572536 484036 577492 484272
rect 572536 477664 572772 484036
rect 573008 477664 573244 484036
rect 573480 477664 573716 484036
rect 573952 477664 574188 484036
rect 574424 477664 574660 484036
rect 574896 477664 575132 484036
rect 575368 477664 575604 484036
rect 575840 477664 576076 484036
rect 576312 477664 576548 484036
rect 576784 477664 577020 484036
rect 577256 477664 577492 484036
rect 562380 455480 567480 455520
rect 562380 455440 562624 455480
rect 562860 455440 563096 455480
rect 563332 455440 563568 455480
rect 563804 455440 564040 455480
rect 564276 455440 564512 455480
rect 564748 455440 564984 455480
rect 565220 455440 565456 455480
rect 565692 455440 565928 455480
rect 566164 455440 566400 455480
rect 566636 455440 566872 455480
rect 567108 455440 567480 455480
rect 562380 455360 562480 455440
rect 562560 455360 562624 455440
rect 562880 455360 562960 455440
rect 563040 455360 563096 455440
rect 563360 455360 563440 455440
rect 563520 455360 563568 455440
rect 563840 455360 563920 455440
rect 564000 455360 564040 455440
rect 564320 455360 564400 455440
rect 564480 455360 564512 455440
rect 564800 455360 564880 455440
rect 564960 455360 564984 455440
rect 565280 455360 565360 455440
rect 565440 455360 565456 455440
rect 565760 455360 565840 455440
rect 565920 455360 565928 455440
rect 566240 455360 566320 455440
rect 566636 455360 566640 455440
rect 566720 455360 566800 455440
rect 567108 455360 567120 455440
rect 567200 455360 567280 455440
rect 567360 455360 567480 455440
rect 562380 455280 562624 455360
rect 562860 455280 563096 455360
rect 563332 455280 563568 455360
rect 563804 455280 564040 455360
rect 564276 455280 564512 455360
rect 564748 455280 564984 455360
rect 565220 455280 565456 455360
rect 565692 455280 565928 455360
rect 566164 455280 566400 455360
rect 566636 455280 566872 455360
rect 567108 455280 567480 455360
rect 562380 455200 562480 455280
rect 562560 455244 562624 455280
rect 562560 455200 562640 455244
rect 562720 455200 562800 455244
rect 562880 455200 562960 455280
rect 563040 455244 563096 455280
rect 563040 455200 563120 455244
rect 563200 455200 563280 455244
rect 563360 455200 563440 455280
rect 563520 455244 563568 455280
rect 563520 455200 563600 455244
rect 563680 455200 563760 455244
rect 563840 455200 563920 455280
rect 564000 455244 564040 455280
rect 564000 455200 564080 455244
rect 564160 455200 564240 455244
rect 564320 455200 564400 455280
rect 564480 455244 564512 455280
rect 564480 455200 564560 455244
rect 564640 455200 564720 455244
rect 564800 455200 564880 455280
rect 564960 455244 564984 455280
rect 564960 455200 565040 455244
rect 565120 455200 565200 455244
rect 565280 455200 565360 455280
rect 565440 455244 565456 455280
rect 565440 455200 565520 455244
rect 565600 455200 565680 455244
rect 565760 455200 565840 455280
rect 565920 455244 565928 455280
rect 565920 455200 566000 455244
rect 566080 455200 566160 455244
rect 566240 455200 566320 455280
rect 566636 455244 566640 455280
rect 566400 455200 566480 455244
rect 566560 455200 566640 455244
rect 566720 455200 566800 455280
rect 567108 455244 567120 455280
rect 566880 455200 566960 455244
rect 567040 455200 567120 455244
rect 567200 455200 567280 455280
rect 567360 455200 567480 455280
rect 562380 455160 567480 455200
rect 572540 455480 577640 455520
rect 572540 455440 572784 455480
rect 573020 455440 573256 455480
rect 573492 455440 573728 455480
rect 573964 455440 574200 455480
rect 574436 455440 574672 455480
rect 574908 455440 575144 455480
rect 575380 455440 575616 455480
rect 575852 455440 576088 455480
rect 576324 455440 576560 455480
rect 576796 455440 577032 455480
rect 577268 455440 577640 455480
rect 572540 455360 572640 455440
rect 572720 455360 572784 455440
rect 573040 455360 573120 455440
rect 573200 455360 573256 455440
rect 573520 455360 573600 455440
rect 573680 455360 573728 455440
rect 574000 455360 574080 455440
rect 574160 455360 574200 455440
rect 574480 455360 574560 455440
rect 574640 455360 574672 455440
rect 574960 455360 575040 455440
rect 575120 455360 575144 455440
rect 575440 455360 575520 455440
rect 575600 455360 575616 455440
rect 575920 455360 576000 455440
rect 576080 455360 576088 455440
rect 576400 455360 576480 455440
rect 576796 455360 576800 455440
rect 576880 455360 576960 455440
rect 577268 455360 577280 455440
rect 577360 455360 577440 455440
rect 577520 455360 577640 455440
rect 572540 455280 572784 455360
rect 573020 455280 573256 455360
rect 573492 455280 573728 455360
rect 573964 455280 574200 455360
rect 574436 455280 574672 455360
rect 574908 455280 575144 455360
rect 575380 455280 575616 455360
rect 575852 455280 576088 455360
rect 576324 455280 576560 455360
rect 576796 455280 577032 455360
rect 577268 455280 577640 455360
rect 572540 455200 572640 455280
rect 572720 455244 572784 455280
rect 572720 455200 572800 455244
rect 572880 455200 572960 455244
rect 573040 455200 573120 455280
rect 573200 455244 573256 455280
rect 573200 455200 573280 455244
rect 573360 455200 573440 455244
rect 573520 455200 573600 455280
rect 573680 455244 573728 455280
rect 573680 455200 573760 455244
rect 573840 455200 573920 455244
rect 574000 455200 574080 455280
rect 574160 455244 574200 455280
rect 574160 455200 574240 455244
rect 574320 455200 574400 455244
rect 574480 455200 574560 455280
rect 574640 455244 574672 455280
rect 574640 455200 574720 455244
rect 574800 455200 574880 455244
rect 574960 455200 575040 455280
rect 575120 455244 575144 455280
rect 575120 455200 575200 455244
rect 575280 455200 575360 455244
rect 575440 455200 575520 455280
rect 575600 455244 575616 455280
rect 575600 455200 575680 455244
rect 575760 455200 575840 455244
rect 575920 455200 576000 455280
rect 576080 455244 576088 455280
rect 576080 455200 576160 455244
rect 576240 455200 576320 455244
rect 576400 455200 576480 455280
rect 576796 455244 576800 455280
rect 576560 455200 576640 455244
rect 576720 455200 576800 455244
rect 576880 455200 576960 455280
rect 577268 455244 577280 455280
rect 577040 455200 577120 455244
rect 577200 455200 577280 455244
rect 577360 455200 577440 455280
rect 577520 455200 577640 455280
rect 572540 455160 577640 455200
rect 572536 426688 577492 426924
rect 572536 420316 572772 426688
rect 573008 420316 573244 426688
rect 573480 420316 573716 426688
rect 573952 420316 574188 426688
rect 574424 420316 574660 426688
rect 574896 420316 575132 426688
rect 575368 420316 575604 426688
rect 575840 420316 576076 426688
rect 576312 420316 576548 426688
rect 576784 420316 577020 426688
rect 577256 420316 577492 426688
rect 477060 377836 483800 378072
rect 477060 377600 477192 377836
rect 477428 377600 477664 377836
rect 477900 377600 478136 377836
rect 478372 377600 478608 377836
rect 478844 377600 479080 377836
rect 479316 377600 479552 377836
rect 479788 377600 480024 377836
rect 480260 377600 480496 377836
rect 480732 377600 480968 377836
rect 481204 377600 481440 377836
rect 481676 377600 481912 377836
rect 482148 377600 482384 377836
rect 482620 377600 482856 377836
rect 483092 377600 483328 377836
rect 483564 377600 483800 377836
rect 477060 377364 483800 377600
rect 477060 377128 477192 377364
rect 477428 377128 477664 377364
rect 477900 377128 478136 377364
rect 478372 377128 478608 377364
rect 478844 377128 479080 377364
rect 479316 377128 479552 377364
rect 479788 377128 480024 377364
rect 480260 377128 480496 377364
rect 480732 377128 480968 377364
rect 481204 377128 481440 377364
rect 481676 377128 481912 377364
rect 482148 377128 482384 377364
rect 482620 377128 482856 377364
rect 483092 377128 483328 377364
rect 483564 377128 483800 377364
rect 477060 376892 483800 377128
rect 477060 376656 477192 376892
rect 477428 376656 477664 376892
rect 477900 376656 478136 376892
rect 478372 376656 478608 376892
rect 478844 376656 479080 376892
rect 479316 376656 479552 376892
rect 479788 376656 480024 376892
rect 480260 376656 480496 376892
rect 480732 376656 480968 376892
rect 481204 376656 481440 376892
rect 481676 376656 481912 376892
rect 482148 376656 482384 376892
rect 482620 376656 482856 376892
rect 483092 376656 483328 376892
rect 483564 376656 483800 376892
rect 477060 376420 483800 376656
rect 477060 376184 477192 376420
rect 477428 376184 477664 376420
rect 477900 376184 478136 376420
rect 478372 376184 478608 376420
rect 478844 376184 479080 376420
rect 479316 376184 479552 376420
rect 479788 376184 480024 376420
rect 480260 376184 480496 376420
rect 480732 376184 480968 376420
rect 481204 376184 481440 376420
rect 481676 376184 481912 376420
rect 482148 376184 482384 376420
rect 482620 376184 482856 376420
rect 483092 376184 483328 376420
rect 483564 376184 483800 376420
rect 477060 375948 483800 376184
rect 477060 375712 477192 375948
rect 477428 375712 477664 375948
rect 477900 375712 478136 375948
rect 478372 375712 478608 375948
rect 478844 375712 479080 375948
rect 479316 375712 479552 375948
rect 479788 375712 480024 375948
rect 480260 375712 480496 375948
rect 480732 375712 480968 375948
rect 481204 375712 481440 375948
rect 481676 375712 481912 375948
rect 482148 375712 482384 375948
rect 482620 375712 482856 375948
rect 483092 375712 483328 375948
rect 483564 375712 483800 375948
rect 477060 375476 483800 375712
rect 477060 375240 477192 375476
rect 477428 375240 477664 375476
rect 477900 375240 478136 375476
rect 478372 375240 478608 375476
rect 478844 375240 479080 375476
rect 479316 375240 479552 375476
rect 479788 375240 480024 375476
rect 480260 375240 480496 375476
rect 480732 375240 480968 375476
rect 481204 375240 481440 375476
rect 481676 375240 481912 375476
rect 482148 375240 482384 375476
rect 482620 375240 482856 375476
rect 483092 375240 483328 375476
rect 483564 375240 483800 375476
rect 477060 375004 483800 375240
rect 477060 374768 477192 375004
rect 477428 374768 477664 375004
rect 477900 374768 478136 375004
rect 478372 374768 478608 375004
rect 478844 374768 479080 375004
rect 479316 374768 479552 375004
rect 479788 374768 480024 375004
rect 480260 374768 480496 375004
rect 480732 374768 480968 375004
rect 481204 374768 481440 375004
rect 481676 374768 481912 375004
rect 482148 374768 482384 375004
rect 482620 374768 482856 375004
rect 483092 374768 483328 375004
rect 483564 374768 483800 375004
rect 477060 374532 483800 374768
rect 477060 374296 477192 374532
rect 477428 374296 477664 374532
rect 477900 374296 478136 374532
rect 478372 374296 478608 374532
rect 478844 374296 479080 374532
rect 479316 374296 479552 374532
rect 479788 374296 480024 374532
rect 480260 374296 480496 374532
rect 480732 374296 480968 374532
rect 481204 374296 481440 374532
rect 481676 374296 481912 374532
rect 482148 374296 482384 374532
rect 482620 374296 482856 374532
rect 483092 374296 483328 374532
rect 483564 374296 483800 374532
rect 477060 374060 483800 374296
rect 477060 373824 477192 374060
rect 477428 373824 477664 374060
rect 477900 373824 478136 374060
rect 478372 373824 478608 374060
rect 478844 373824 479080 374060
rect 479316 373824 479552 374060
rect 479788 373824 480024 374060
rect 480260 373824 480496 374060
rect 480732 373824 480968 374060
rect 481204 373824 481440 374060
rect 481676 373824 481912 374060
rect 482148 373824 482384 374060
rect 482620 373824 482856 374060
rect 483092 373824 483328 374060
rect 483564 373824 483800 374060
rect 477060 373588 483800 373824
rect 477060 373352 477192 373588
rect 477428 373352 477664 373588
rect 477900 373352 478136 373588
rect 478372 373352 478608 373588
rect 478844 373352 479080 373588
rect 479316 373352 479552 373588
rect 479788 373352 480024 373588
rect 480260 373352 480496 373588
rect 480732 373352 480968 373588
rect 481204 373352 481440 373588
rect 481676 373352 481912 373588
rect 482148 373352 482384 373588
rect 482620 373352 482856 373588
rect 483092 373352 483328 373588
rect 483564 373352 483800 373588
rect 477060 373116 483800 373352
rect 477060 372880 477192 373116
rect 477428 372880 477664 373116
rect 477900 372880 478136 373116
rect 478372 372880 478608 373116
rect 478844 372880 479080 373116
rect 479316 372880 479552 373116
rect 479788 372880 480024 373116
rect 480260 372880 480496 373116
rect 480732 372880 480968 373116
rect 481204 372880 481440 373116
rect 481676 372880 481912 373116
rect 482148 372880 482384 373116
rect 482620 372880 482856 373116
rect 483092 372880 483328 373116
rect 483564 372880 483800 373116
rect 477060 372644 483800 372880
rect 477060 372408 477192 372644
rect 477428 372408 477664 372644
rect 477900 372408 478136 372644
rect 478372 372408 478608 372644
rect 478844 372408 479080 372644
rect 479316 372408 479552 372644
rect 479788 372408 480024 372644
rect 480260 372408 480496 372644
rect 480732 372408 480968 372644
rect 481204 372408 481440 372644
rect 481676 372408 481912 372644
rect 482148 372408 482384 372644
rect 482620 372408 482856 372644
rect 483092 372408 483328 372644
rect 483564 372408 483800 372644
rect 477060 372172 483800 372408
rect 477060 371936 477192 372172
rect 477428 371936 477664 372172
rect 477900 371936 478136 372172
rect 478372 371936 478608 372172
rect 478844 371936 479080 372172
rect 479316 371936 479552 372172
rect 479788 371936 480024 372172
rect 480260 371936 480496 372172
rect 480732 371936 480968 372172
rect 481204 371936 481440 372172
rect 481676 371936 481912 372172
rect 482148 371936 482384 372172
rect 482620 371936 482856 372172
rect 483092 371936 483328 372172
rect 483564 371936 483800 372172
rect 477060 371700 483800 371936
rect 477060 371464 477192 371700
rect 477428 371464 477664 371700
rect 477900 371464 478136 371700
rect 478372 371464 478608 371700
rect 478844 371464 479080 371700
rect 479316 371464 479552 371700
rect 479788 371464 480024 371700
rect 480260 371464 480496 371700
rect 480732 371464 480968 371700
rect 481204 371464 481440 371700
rect 481676 371464 481912 371700
rect 482148 371464 482384 371700
rect 482620 371464 482856 371700
rect 483092 371464 483328 371700
rect 483564 371464 483800 371700
rect 562388 377600 567816 378072
rect 477060 371200 483726 371464
rect 562388 371228 562624 377600
rect 562860 371228 563096 377600
rect 563332 371228 563568 377600
rect 563804 371228 564040 377600
rect 564276 371228 564512 377600
rect 564748 371228 564984 377600
rect 565220 371228 565456 377600
rect 565692 371228 565928 377600
rect 566164 371228 566400 377600
rect 566636 371228 566872 377600
rect 567108 371228 567816 377600
rect 562388 370992 567816 371228
<< via4 >>
rect 572772 696908 573008 697144
rect 573244 696908 573480 697144
rect 573716 696908 573952 697144
rect 574188 696908 574424 697144
rect 574660 696908 574896 697144
rect 575132 696908 575368 697144
rect 575604 696908 575840 697144
rect 576076 696908 576312 697144
rect 576548 696908 576784 697144
rect 577020 696908 577256 697144
rect 572772 696436 573008 696672
rect 573244 696436 573480 696672
rect 573716 696436 573952 696672
rect 574188 696436 574424 696672
rect 574660 696436 574896 696672
rect 575132 696436 575368 696672
rect 575604 696436 575840 696672
rect 576076 696436 576312 696672
rect 576548 696436 576784 696672
rect 577020 696436 577256 696672
rect 572772 695964 573008 696200
rect 573244 695964 573480 696200
rect 573716 695964 573952 696200
rect 574188 695964 574424 696200
rect 574660 695964 574896 696200
rect 575132 695964 575368 696200
rect 575604 695964 575840 696200
rect 576076 695964 576312 696200
rect 576548 695964 576784 696200
rect 577020 695964 577256 696200
rect 572772 695492 573008 695728
rect 573244 695492 573480 695728
rect 573716 695492 573952 695728
rect 574188 695492 574424 695728
rect 574660 695492 574896 695728
rect 575132 695492 575368 695728
rect 575604 695492 575840 695728
rect 576076 695492 576312 695728
rect 576548 695492 576784 695728
rect 577020 695492 577256 695728
rect 572772 695020 573008 695256
rect 573244 695020 573480 695256
rect 573716 695020 573952 695256
rect 574188 695020 574424 695256
rect 574660 695020 574896 695256
rect 575132 695020 575368 695256
rect 575604 695020 575840 695256
rect 576076 695020 576312 695256
rect 576548 695020 576784 695256
rect 577020 695020 577256 695256
rect 572772 694548 573008 694784
rect 573244 694548 573480 694784
rect 573716 694548 573952 694784
rect 574188 694548 574424 694784
rect 574660 694548 574896 694784
rect 575132 694548 575368 694784
rect 575604 694548 575840 694784
rect 576076 694548 576312 694784
rect 576548 694548 576784 694784
rect 577020 694548 577256 694784
rect 572772 694076 573008 694312
rect 573244 694076 573480 694312
rect 573716 694076 573952 694312
rect 574188 694076 574424 694312
rect 574660 694076 574896 694312
rect 575132 694076 575368 694312
rect 575604 694076 575840 694312
rect 576076 694076 576312 694312
rect 576548 694076 576784 694312
rect 577020 694076 577256 694312
rect 572772 693604 573008 693840
rect 573244 693604 573480 693840
rect 573716 693604 573952 693840
rect 574188 693604 574424 693840
rect 574660 693604 574896 693840
rect 575132 693604 575368 693840
rect 575604 693604 575840 693840
rect 576076 693604 576312 693840
rect 576548 693604 576784 693840
rect 577020 693604 577256 693840
rect 572772 693132 573008 693368
rect 573244 693132 573480 693368
rect 573716 693132 573952 693368
rect 574188 693132 574424 693368
rect 574660 693132 574896 693368
rect 575132 693132 575368 693368
rect 575604 693132 575840 693368
rect 576076 693132 576312 693368
rect 576548 693132 576784 693368
rect 577020 693132 577256 693368
rect 572772 692660 573008 692896
rect 573244 692660 573480 692896
rect 573716 692660 573952 692896
rect 574188 692660 574424 692896
rect 574660 692660 574896 692896
rect 575132 692660 575368 692896
rect 575604 692660 575840 692896
rect 576076 692660 576312 692896
rect 576548 692660 576784 692896
rect 577020 692660 577256 692896
rect 562480 644524 567400 644584
rect 562480 639844 562600 644524
rect 562600 639844 567400 644524
rect 562480 639784 567400 639844
rect 562480 634524 567400 634584
rect 562480 629844 562600 634524
rect 562600 629844 567400 634524
rect 562480 629784 567400 629844
rect 562624 522268 562860 522504
rect 562624 521796 562860 522032
rect 562624 521324 562860 521560
rect 562624 520852 562860 521088
rect 562624 520380 562860 520616
rect 562624 519908 562860 520144
rect 562624 519436 562860 519672
rect 562624 518964 562860 519200
rect 562624 518492 562860 518728
rect 562624 518020 562860 518256
rect 562624 517548 562860 517784
rect 562624 517076 562860 517312
rect 562624 516604 562860 516840
rect 563096 522268 563332 522504
rect 563096 521796 563332 522032
rect 563096 521324 563332 521560
rect 563096 520852 563332 521088
rect 563096 520380 563332 520616
rect 563096 519908 563332 520144
rect 563096 519436 563332 519672
rect 563096 518964 563332 519200
rect 563096 518492 563332 518728
rect 563096 518020 563332 518256
rect 563096 517548 563332 517784
rect 563096 517076 563332 517312
rect 563096 516604 563332 516840
rect 563568 522268 563804 522504
rect 563568 521796 563804 522032
rect 563568 521324 563804 521560
rect 563568 520852 563804 521088
rect 563568 520380 563804 520616
rect 563568 519908 563804 520144
rect 563568 519436 563804 519672
rect 563568 518964 563804 519200
rect 563568 518492 563804 518728
rect 563568 518020 563804 518256
rect 563568 517548 563804 517784
rect 563568 517076 563804 517312
rect 563568 516604 563804 516840
rect 564040 522268 564276 522504
rect 564040 521796 564276 522032
rect 564040 521324 564276 521560
rect 564040 520852 564276 521088
rect 564040 520380 564276 520616
rect 564040 519908 564276 520144
rect 564040 519436 564276 519672
rect 564040 518964 564276 519200
rect 564040 518492 564276 518728
rect 564040 518020 564276 518256
rect 564040 517548 564276 517784
rect 564040 517076 564276 517312
rect 564040 516604 564276 516840
rect 564512 522268 564748 522504
rect 564512 521796 564748 522032
rect 564512 521324 564748 521560
rect 564512 520852 564748 521088
rect 564512 520380 564748 520616
rect 564512 519908 564748 520144
rect 564512 519436 564748 519672
rect 564512 518964 564748 519200
rect 564512 518492 564748 518728
rect 564512 518020 564748 518256
rect 564512 517548 564748 517784
rect 564512 517076 564748 517312
rect 564512 516604 564748 516840
rect 564984 522268 565220 522504
rect 564984 521796 565220 522032
rect 564984 521324 565220 521560
rect 564984 520852 565220 521088
rect 564984 520380 565220 520616
rect 564984 519908 565220 520144
rect 564984 519436 565220 519672
rect 564984 518964 565220 519200
rect 564984 518492 565220 518728
rect 564984 518020 565220 518256
rect 564984 517548 565220 517784
rect 564984 517076 565220 517312
rect 564984 516604 565220 516840
rect 565456 522268 565692 522504
rect 565456 521796 565692 522032
rect 565456 521324 565692 521560
rect 565456 520852 565692 521088
rect 565456 520380 565692 520616
rect 565456 519908 565692 520144
rect 565456 519436 565692 519672
rect 565456 518964 565692 519200
rect 565456 518492 565692 518728
rect 565456 518020 565692 518256
rect 565456 517548 565692 517784
rect 565456 517076 565692 517312
rect 565456 516604 565692 516840
rect 565928 522268 566164 522504
rect 565928 521796 566164 522032
rect 565928 521324 566164 521560
rect 565928 520852 566164 521088
rect 565928 520380 566164 520616
rect 565928 519908 566164 520144
rect 565928 519436 566164 519672
rect 565928 518964 566164 519200
rect 565928 518492 566164 518728
rect 565928 518020 566164 518256
rect 565928 517548 566164 517784
rect 565928 517076 566164 517312
rect 565928 516604 566164 516840
rect 566400 522268 566636 522504
rect 566400 521796 566636 522032
rect 566400 521324 566636 521560
rect 566400 520852 566636 521088
rect 566400 520380 566636 520616
rect 566400 519908 566636 520144
rect 566400 519436 566636 519672
rect 566400 518964 566636 519200
rect 566400 518492 566636 518728
rect 566400 518020 566636 518256
rect 566400 517548 566636 517784
rect 566400 517076 566636 517312
rect 566400 516604 566636 516840
rect 566872 522268 567108 522504
rect 566872 521796 567108 522032
rect 566872 521324 567108 521560
rect 566872 520852 567108 521088
rect 566872 520380 567108 520616
rect 566872 519908 567108 520144
rect 566872 519436 567108 519672
rect 566872 518964 567108 519200
rect 566872 518492 567108 518728
rect 566872 518020 567108 518256
rect 566872 517548 567108 517784
rect 566872 517076 567108 517312
rect 566872 516604 567108 516840
rect 562624 495742 562860 495782
rect 563096 495742 563332 495782
rect 563568 495742 563804 495782
rect 564040 495742 564276 495782
rect 564512 495742 564748 495782
rect 564984 495742 565220 495782
rect 565456 495742 565692 495782
rect 565928 495742 566164 495782
rect 566400 495742 566636 495782
rect 566872 495742 567108 495782
rect 562624 495662 562640 495742
rect 562640 495662 562720 495742
rect 562720 495662 562800 495742
rect 562800 495662 562860 495742
rect 563096 495662 563120 495742
rect 563120 495662 563200 495742
rect 563200 495662 563280 495742
rect 563280 495662 563332 495742
rect 563568 495662 563600 495742
rect 563600 495662 563680 495742
rect 563680 495662 563760 495742
rect 563760 495662 563804 495742
rect 564040 495662 564080 495742
rect 564080 495662 564160 495742
rect 564160 495662 564240 495742
rect 564240 495662 564276 495742
rect 564512 495662 564560 495742
rect 564560 495662 564640 495742
rect 564640 495662 564720 495742
rect 564720 495662 564748 495742
rect 564984 495662 565040 495742
rect 565040 495662 565120 495742
rect 565120 495662 565200 495742
rect 565200 495662 565220 495742
rect 565456 495662 565520 495742
rect 565520 495662 565600 495742
rect 565600 495662 565680 495742
rect 565680 495662 565692 495742
rect 565928 495662 566000 495742
rect 566000 495662 566080 495742
rect 566080 495662 566160 495742
rect 566160 495662 566164 495742
rect 566400 495662 566480 495742
rect 566480 495662 566560 495742
rect 566560 495662 566636 495742
rect 566872 495662 566880 495742
rect 566880 495662 566960 495742
rect 566960 495662 567040 495742
rect 567040 495662 567108 495742
rect 562624 495582 562860 495662
rect 563096 495582 563332 495662
rect 563568 495582 563804 495662
rect 564040 495582 564276 495662
rect 564512 495582 564748 495662
rect 564984 495582 565220 495662
rect 565456 495582 565692 495662
rect 565928 495582 566164 495662
rect 566400 495582 566636 495662
rect 566872 495582 567108 495662
rect 562624 495546 562640 495582
rect 562640 495546 562720 495582
rect 562720 495546 562800 495582
rect 562800 495546 562860 495582
rect 563096 495546 563120 495582
rect 563120 495546 563200 495582
rect 563200 495546 563280 495582
rect 563280 495546 563332 495582
rect 563568 495546 563600 495582
rect 563600 495546 563680 495582
rect 563680 495546 563760 495582
rect 563760 495546 563804 495582
rect 564040 495546 564080 495582
rect 564080 495546 564160 495582
rect 564160 495546 564240 495582
rect 564240 495546 564276 495582
rect 564512 495546 564560 495582
rect 564560 495546 564640 495582
rect 564640 495546 564720 495582
rect 564720 495546 564748 495582
rect 564984 495546 565040 495582
rect 565040 495546 565120 495582
rect 565120 495546 565200 495582
rect 565200 495546 565220 495582
rect 565456 495546 565520 495582
rect 565520 495546 565600 495582
rect 565600 495546 565680 495582
rect 565680 495546 565692 495582
rect 565928 495546 566000 495582
rect 566000 495546 566080 495582
rect 566080 495546 566160 495582
rect 566160 495546 566164 495582
rect 566400 495546 566480 495582
rect 566480 495546 566560 495582
rect 566560 495546 566636 495582
rect 566872 495546 566880 495582
rect 566880 495546 566960 495582
rect 566960 495546 567040 495582
rect 567040 495546 567108 495582
rect 572784 495742 573020 495782
rect 573256 495742 573492 495782
rect 573728 495742 573964 495782
rect 574200 495742 574436 495782
rect 574672 495742 574908 495782
rect 575144 495742 575380 495782
rect 575616 495742 575852 495782
rect 576088 495742 576324 495782
rect 576560 495742 576796 495782
rect 577032 495742 577268 495782
rect 572784 495662 572800 495742
rect 572800 495662 572880 495742
rect 572880 495662 572960 495742
rect 572960 495662 573020 495742
rect 573256 495662 573280 495742
rect 573280 495662 573360 495742
rect 573360 495662 573440 495742
rect 573440 495662 573492 495742
rect 573728 495662 573760 495742
rect 573760 495662 573840 495742
rect 573840 495662 573920 495742
rect 573920 495662 573964 495742
rect 574200 495662 574240 495742
rect 574240 495662 574320 495742
rect 574320 495662 574400 495742
rect 574400 495662 574436 495742
rect 574672 495662 574720 495742
rect 574720 495662 574800 495742
rect 574800 495662 574880 495742
rect 574880 495662 574908 495742
rect 575144 495662 575200 495742
rect 575200 495662 575280 495742
rect 575280 495662 575360 495742
rect 575360 495662 575380 495742
rect 575616 495662 575680 495742
rect 575680 495662 575760 495742
rect 575760 495662 575840 495742
rect 575840 495662 575852 495742
rect 576088 495662 576160 495742
rect 576160 495662 576240 495742
rect 576240 495662 576320 495742
rect 576320 495662 576324 495742
rect 576560 495662 576640 495742
rect 576640 495662 576720 495742
rect 576720 495662 576796 495742
rect 577032 495662 577040 495742
rect 577040 495662 577120 495742
rect 577120 495662 577200 495742
rect 577200 495662 577268 495742
rect 572784 495582 573020 495662
rect 573256 495582 573492 495662
rect 573728 495582 573964 495662
rect 574200 495582 574436 495662
rect 574672 495582 574908 495662
rect 575144 495582 575380 495662
rect 575616 495582 575852 495662
rect 576088 495582 576324 495662
rect 576560 495582 576796 495662
rect 577032 495582 577268 495662
rect 572784 495546 572800 495582
rect 572800 495546 572880 495582
rect 572880 495546 572960 495582
rect 572960 495546 573020 495582
rect 573256 495546 573280 495582
rect 573280 495546 573360 495582
rect 573360 495546 573440 495582
rect 573440 495546 573492 495582
rect 573728 495546 573760 495582
rect 573760 495546 573840 495582
rect 573840 495546 573920 495582
rect 573920 495546 573964 495582
rect 574200 495546 574240 495582
rect 574240 495546 574320 495582
rect 574320 495546 574400 495582
rect 574400 495546 574436 495582
rect 574672 495546 574720 495582
rect 574720 495546 574800 495582
rect 574800 495546 574880 495582
rect 574880 495546 574908 495582
rect 575144 495546 575200 495582
rect 575200 495546 575280 495582
rect 575280 495546 575360 495582
rect 575360 495546 575380 495582
rect 575616 495546 575680 495582
rect 575680 495546 575760 495582
rect 575760 495546 575840 495582
rect 575840 495546 575852 495582
rect 576088 495546 576160 495582
rect 576160 495546 576240 495582
rect 576240 495546 576320 495582
rect 576320 495546 576324 495582
rect 576560 495546 576640 495582
rect 576640 495546 576720 495582
rect 576720 495546 576796 495582
rect 577032 495546 577040 495582
rect 577040 495546 577120 495582
rect 577120 495546 577200 495582
rect 577200 495546 577268 495582
rect 572772 483800 573008 484036
rect 572772 483328 573008 483564
rect 572772 482856 573008 483092
rect 572772 482384 573008 482620
rect 572772 481912 573008 482148
rect 572772 481440 573008 481676
rect 572772 480968 573008 481204
rect 572772 480496 573008 480732
rect 572772 480024 573008 480260
rect 572772 479552 573008 479788
rect 572772 479080 573008 479316
rect 572772 478608 573008 478844
rect 572772 478136 573008 478372
rect 572772 477664 573008 477900
rect 573244 483800 573480 484036
rect 573244 483328 573480 483564
rect 573244 482856 573480 483092
rect 573244 482384 573480 482620
rect 573244 481912 573480 482148
rect 573244 481440 573480 481676
rect 573244 480968 573480 481204
rect 573244 480496 573480 480732
rect 573244 480024 573480 480260
rect 573244 479552 573480 479788
rect 573244 479080 573480 479316
rect 573244 478608 573480 478844
rect 573244 478136 573480 478372
rect 573244 477664 573480 477900
rect 573716 483800 573952 484036
rect 573716 483328 573952 483564
rect 573716 482856 573952 483092
rect 573716 482384 573952 482620
rect 573716 481912 573952 482148
rect 573716 481440 573952 481676
rect 573716 480968 573952 481204
rect 573716 480496 573952 480732
rect 573716 480024 573952 480260
rect 573716 479552 573952 479788
rect 573716 479080 573952 479316
rect 573716 478608 573952 478844
rect 573716 478136 573952 478372
rect 573716 477664 573952 477900
rect 574188 483800 574424 484036
rect 574188 483328 574424 483564
rect 574188 482856 574424 483092
rect 574188 482384 574424 482620
rect 574188 481912 574424 482148
rect 574188 481440 574424 481676
rect 574188 480968 574424 481204
rect 574188 480496 574424 480732
rect 574188 480024 574424 480260
rect 574188 479552 574424 479788
rect 574188 479080 574424 479316
rect 574188 478608 574424 478844
rect 574188 478136 574424 478372
rect 574188 477664 574424 477900
rect 574660 483800 574896 484036
rect 574660 483328 574896 483564
rect 574660 482856 574896 483092
rect 574660 482384 574896 482620
rect 574660 481912 574896 482148
rect 574660 481440 574896 481676
rect 574660 480968 574896 481204
rect 574660 480496 574896 480732
rect 574660 480024 574896 480260
rect 574660 479552 574896 479788
rect 574660 479080 574896 479316
rect 574660 478608 574896 478844
rect 574660 478136 574896 478372
rect 574660 477664 574896 477900
rect 575132 483800 575368 484036
rect 575132 483328 575368 483564
rect 575132 482856 575368 483092
rect 575132 482384 575368 482620
rect 575132 481912 575368 482148
rect 575132 481440 575368 481676
rect 575132 480968 575368 481204
rect 575132 480496 575368 480732
rect 575132 480024 575368 480260
rect 575132 479552 575368 479788
rect 575132 479080 575368 479316
rect 575132 478608 575368 478844
rect 575132 478136 575368 478372
rect 575132 477664 575368 477900
rect 575604 483800 575840 484036
rect 575604 483328 575840 483564
rect 575604 482856 575840 483092
rect 575604 482384 575840 482620
rect 575604 481912 575840 482148
rect 575604 481440 575840 481676
rect 575604 480968 575840 481204
rect 575604 480496 575840 480732
rect 575604 480024 575840 480260
rect 575604 479552 575840 479788
rect 575604 479080 575840 479316
rect 575604 478608 575840 478844
rect 575604 478136 575840 478372
rect 575604 477664 575840 477900
rect 576076 483800 576312 484036
rect 576076 483328 576312 483564
rect 576076 482856 576312 483092
rect 576076 482384 576312 482620
rect 576076 481912 576312 482148
rect 576076 481440 576312 481676
rect 576076 480968 576312 481204
rect 576076 480496 576312 480732
rect 576076 480024 576312 480260
rect 576076 479552 576312 479788
rect 576076 479080 576312 479316
rect 576076 478608 576312 478844
rect 576076 478136 576312 478372
rect 576076 477664 576312 477900
rect 576548 483800 576784 484036
rect 576548 483328 576784 483564
rect 576548 482856 576784 483092
rect 576548 482384 576784 482620
rect 576548 481912 576784 482148
rect 576548 481440 576784 481676
rect 576548 480968 576784 481204
rect 576548 480496 576784 480732
rect 576548 480024 576784 480260
rect 576548 479552 576784 479788
rect 576548 479080 576784 479316
rect 576548 478608 576784 478844
rect 576548 478136 576784 478372
rect 576548 477664 576784 477900
rect 577020 483800 577256 484036
rect 577020 483328 577256 483564
rect 577020 482856 577256 483092
rect 577020 482384 577256 482620
rect 577020 481912 577256 482148
rect 577020 481440 577256 481676
rect 577020 480968 577256 481204
rect 577020 480496 577256 480732
rect 577020 480024 577256 480260
rect 577020 479552 577256 479788
rect 577020 479080 577256 479316
rect 577020 478608 577256 478844
rect 577020 478136 577256 478372
rect 577020 477664 577256 477900
rect 562624 455440 562860 455480
rect 563096 455440 563332 455480
rect 563568 455440 563804 455480
rect 564040 455440 564276 455480
rect 564512 455440 564748 455480
rect 564984 455440 565220 455480
rect 565456 455440 565692 455480
rect 565928 455440 566164 455480
rect 566400 455440 566636 455480
rect 566872 455440 567108 455480
rect 562624 455360 562640 455440
rect 562640 455360 562720 455440
rect 562720 455360 562800 455440
rect 562800 455360 562860 455440
rect 563096 455360 563120 455440
rect 563120 455360 563200 455440
rect 563200 455360 563280 455440
rect 563280 455360 563332 455440
rect 563568 455360 563600 455440
rect 563600 455360 563680 455440
rect 563680 455360 563760 455440
rect 563760 455360 563804 455440
rect 564040 455360 564080 455440
rect 564080 455360 564160 455440
rect 564160 455360 564240 455440
rect 564240 455360 564276 455440
rect 564512 455360 564560 455440
rect 564560 455360 564640 455440
rect 564640 455360 564720 455440
rect 564720 455360 564748 455440
rect 564984 455360 565040 455440
rect 565040 455360 565120 455440
rect 565120 455360 565200 455440
rect 565200 455360 565220 455440
rect 565456 455360 565520 455440
rect 565520 455360 565600 455440
rect 565600 455360 565680 455440
rect 565680 455360 565692 455440
rect 565928 455360 566000 455440
rect 566000 455360 566080 455440
rect 566080 455360 566160 455440
rect 566160 455360 566164 455440
rect 566400 455360 566480 455440
rect 566480 455360 566560 455440
rect 566560 455360 566636 455440
rect 566872 455360 566880 455440
rect 566880 455360 566960 455440
rect 566960 455360 567040 455440
rect 567040 455360 567108 455440
rect 562624 455280 562860 455360
rect 563096 455280 563332 455360
rect 563568 455280 563804 455360
rect 564040 455280 564276 455360
rect 564512 455280 564748 455360
rect 564984 455280 565220 455360
rect 565456 455280 565692 455360
rect 565928 455280 566164 455360
rect 566400 455280 566636 455360
rect 566872 455280 567108 455360
rect 562624 455244 562640 455280
rect 562640 455244 562720 455280
rect 562720 455244 562800 455280
rect 562800 455244 562860 455280
rect 563096 455244 563120 455280
rect 563120 455244 563200 455280
rect 563200 455244 563280 455280
rect 563280 455244 563332 455280
rect 563568 455244 563600 455280
rect 563600 455244 563680 455280
rect 563680 455244 563760 455280
rect 563760 455244 563804 455280
rect 564040 455244 564080 455280
rect 564080 455244 564160 455280
rect 564160 455244 564240 455280
rect 564240 455244 564276 455280
rect 564512 455244 564560 455280
rect 564560 455244 564640 455280
rect 564640 455244 564720 455280
rect 564720 455244 564748 455280
rect 564984 455244 565040 455280
rect 565040 455244 565120 455280
rect 565120 455244 565200 455280
rect 565200 455244 565220 455280
rect 565456 455244 565520 455280
rect 565520 455244 565600 455280
rect 565600 455244 565680 455280
rect 565680 455244 565692 455280
rect 565928 455244 566000 455280
rect 566000 455244 566080 455280
rect 566080 455244 566160 455280
rect 566160 455244 566164 455280
rect 566400 455244 566480 455280
rect 566480 455244 566560 455280
rect 566560 455244 566636 455280
rect 566872 455244 566880 455280
rect 566880 455244 566960 455280
rect 566960 455244 567040 455280
rect 567040 455244 567108 455280
rect 572784 455440 573020 455480
rect 573256 455440 573492 455480
rect 573728 455440 573964 455480
rect 574200 455440 574436 455480
rect 574672 455440 574908 455480
rect 575144 455440 575380 455480
rect 575616 455440 575852 455480
rect 576088 455440 576324 455480
rect 576560 455440 576796 455480
rect 577032 455440 577268 455480
rect 572784 455360 572800 455440
rect 572800 455360 572880 455440
rect 572880 455360 572960 455440
rect 572960 455360 573020 455440
rect 573256 455360 573280 455440
rect 573280 455360 573360 455440
rect 573360 455360 573440 455440
rect 573440 455360 573492 455440
rect 573728 455360 573760 455440
rect 573760 455360 573840 455440
rect 573840 455360 573920 455440
rect 573920 455360 573964 455440
rect 574200 455360 574240 455440
rect 574240 455360 574320 455440
rect 574320 455360 574400 455440
rect 574400 455360 574436 455440
rect 574672 455360 574720 455440
rect 574720 455360 574800 455440
rect 574800 455360 574880 455440
rect 574880 455360 574908 455440
rect 575144 455360 575200 455440
rect 575200 455360 575280 455440
rect 575280 455360 575360 455440
rect 575360 455360 575380 455440
rect 575616 455360 575680 455440
rect 575680 455360 575760 455440
rect 575760 455360 575840 455440
rect 575840 455360 575852 455440
rect 576088 455360 576160 455440
rect 576160 455360 576240 455440
rect 576240 455360 576320 455440
rect 576320 455360 576324 455440
rect 576560 455360 576640 455440
rect 576640 455360 576720 455440
rect 576720 455360 576796 455440
rect 577032 455360 577040 455440
rect 577040 455360 577120 455440
rect 577120 455360 577200 455440
rect 577200 455360 577268 455440
rect 572784 455280 573020 455360
rect 573256 455280 573492 455360
rect 573728 455280 573964 455360
rect 574200 455280 574436 455360
rect 574672 455280 574908 455360
rect 575144 455280 575380 455360
rect 575616 455280 575852 455360
rect 576088 455280 576324 455360
rect 576560 455280 576796 455360
rect 577032 455280 577268 455360
rect 572784 455244 572800 455280
rect 572800 455244 572880 455280
rect 572880 455244 572960 455280
rect 572960 455244 573020 455280
rect 573256 455244 573280 455280
rect 573280 455244 573360 455280
rect 573360 455244 573440 455280
rect 573440 455244 573492 455280
rect 573728 455244 573760 455280
rect 573760 455244 573840 455280
rect 573840 455244 573920 455280
rect 573920 455244 573964 455280
rect 574200 455244 574240 455280
rect 574240 455244 574320 455280
rect 574320 455244 574400 455280
rect 574400 455244 574436 455280
rect 574672 455244 574720 455280
rect 574720 455244 574800 455280
rect 574800 455244 574880 455280
rect 574880 455244 574908 455280
rect 575144 455244 575200 455280
rect 575200 455244 575280 455280
rect 575280 455244 575360 455280
rect 575360 455244 575380 455280
rect 575616 455244 575680 455280
rect 575680 455244 575760 455280
rect 575760 455244 575840 455280
rect 575840 455244 575852 455280
rect 576088 455244 576160 455280
rect 576160 455244 576240 455280
rect 576240 455244 576320 455280
rect 576320 455244 576324 455280
rect 576560 455244 576640 455280
rect 576640 455244 576720 455280
rect 576720 455244 576796 455280
rect 577032 455244 577040 455280
rect 577040 455244 577120 455280
rect 577120 455244 577200 455280
rect 577200 455244 577268 455280
rect 572772 426452 573008 426688
rect 572772 425980 573008 426216
rect 572772 425508 573008 425744
rect 572772 425036 573008 425272
rect 572772 424564 573008 424800
rect 572772 424092 573008 424328
rect 572772 423620 573008 423856
rect 572772 423148 573008 423384
rect 572772 422676 573008 422912
rect 572772 422204 573008 422440
rect 572772 421732 573008 421968
rect 572772 421260 573008 421496
rect 572772 420788 573008 421024
rect 572772 420316 573008 420552
rect 573244 426452 573480 426688
rect 573244 425980 573480 426216
rect 573244 425508 573480 425744
rect 573244 425036 573480 425272
rect 573244 424564 573480 424800
rect 573244 424092 573480 424328
rect 573244 423620 573480 423856
rect 573244 423148 573480 423384
rect 573244 422676 573480 422912
rect 573244 422204 573480 422440
rect 573244 421732 573480 421968
rect 573244 421260 573480 421496
rect 573244 420788 573480 421024
rect 573244 420316 573480 420552
rect 573716 426452 573952 426688
rect 573716 425980 573952 426216
rect 573716 425508 573952 425744
rect 573716 425036 573952 425272
rect 573716 424564 573952 424800
rect 573716 424092 573952 424328
rect 573716 423620 573952 423856
rect 573716 423148 573952 423384
rect 573716 422676 573952 422912
rect 573716 422204 573952 422440
rect 573716 421732 573952 421968
rect 573716 421260 573952 421496
rect 573716 420788 573952 421024
rect 573716 420316 573952 420552
rect 574188 426452 574424 426688
rect 574188 425980 574424 426216
rect 574188 425508 574424 425744
rect 574188 425036 574424 425272
rect 574188 424564 574424 424800
rect 574188 424092 574424 424328
rect 574188 423620 574424 423856
rect 574188 423148 574424 423384
rect 574188 422676 574424 422912
rect 574188 422204 574424 422440
rect 574188 421732 574424 421968
rect 574188 421260 574424 421496
rect 574188 420788 574424 421024
rect 574188 420316 574424 420552
rect 574660 426452 574896 426688
rect 574660 425980 574896 426216
rect 574660 425508 574896 425744
rect 574660 425036 574896 425272
rect 574660 424564 574896 424800
rect 574660 424092 574896 424328
rect 574660 423620 574896 423856
rect 574660 423148 574896 423384
rect 574660 422676 574896 422912
rect 574660 422204 574896 422440
rect 574660 421732 574896 421968
rect 574660 421260 574896 421496
rect 574660 420788 574896 421024
rect 574660 420316 574896 420552
rect 575132 426452 575368 426688
rect 575132 425980 575368 426216
rect 575132 425508 575368 425744
rect 575132 425036 575368 425272
rect 575132 424564 575368 424800
rect 575132 424092 575368 424328
rect 575132 423620 575368 423856
rect 575132 423148 575368 423384
rect 575132 422676 575368 422912
rect 575132 422204 575368 422440
rect 575132 421732 575368 421968
rect 575132 421260 575368 421496
rect 575132 420788 575368 421024
rect 575132 420316 575368 420552
rect 575604 426452 575840 426688
rect 575604 425980 575840 426216
rect 575604 425508 575840 425744
rect 575604 425036 575840 425272
rect 575604 424564 575840 424800
rect 575604 424092 575840 424328
rect 575604 423620 575840 423856
rect 575604 423148 575840 423384
rect 575604 422676 575840 422912
rect 575604 422204 575840 422440
rect 575604 421732 575840 421968
rect 575604 421260 575840 421496
rect 575604 420788 575840 421024
rect 575604 420316 575840 420552
rect 576076 426452 576312 426688
rect 576076 425980 576312 426216
rect 576076 425508 576312 425744
rect 576076 425036 576312 425272
rect 576076 424564 576312 424800
rect 576076 424092 576312 424328
rect 576076 423620 576312 423856
rect 576076 423148 576312 423384
rect 576076 422676 576312 422912
rect 576076 422204 576312 422440
rect 576076 421732 576312 421968
rect 576076 421260 576312 421496
rect 576076 420788 576312 421024
rect 576076 420316 576312 420552
rect 576548 426452 576784 426688
rect 576548 425980 576784 426216
rect 576548 425508 576784 425744
rect 576548 425036 576784 425272
rect 576548 424564 576784 424800
rect 576548 424092 576784 424328
rect 576548 423620 576784 423856
rect 576548 423148 576784 423384
rect 576548 422676 576784 422912
rect 576548 422204 576784 422440
rect 576548 421732 576784 421968
rect 576548 421260 576784 421496
rect 576548 420788 576784 421024
rect 576548 420316 576784 420552
rect 577020 426452 577256 426688
rect 577020 425980 577256 426216
rect 577020 425508 577256 425744
rect 577020 425036 577256 425272
rect 577020 424564 577256 424800
rect 577020 424092 577256 424328
rect 577020 423620 577256 423856
rect 577020 423148 577256 423384
rect 577020 422676 577256 422912
rect 577020 422204 577256 422440
rect 577020 421732 577256 421968
rect 577020 421260 577256 421496
rect 577020 420788 577256 421024
rect 577020 420316 577256 420552
rect 562624 377128 562860 377364
rect 562624 376656 562860 376892
rect 562624 376184 562860 376420
rect 562624 375712 562860 375948
rect 562624 375240 562860 375476
rect 562624 374768 562860 375004
rect 562624 374296 562860 374532
rect 562624 373824 562860 374060
rect 562624 373352 562860 373588
rect 562624 372880 562860 373116
rect 562624 372408 562860 372644
rect 562624 371936 562860 372172
rect 562624 371464 562860 371700
rect 563096 377128 563332 377364
rect 563096 376656 563332 376892
rect 563096 376184 563332 376420
rect 563096 375712 563332 375948
rect 563096 375240 563332 375476
rect 563096 374768 563332 375004
rect 563096 374296 563332 374532
rect 563096 373824 563332 374060
rect 563096 373352 563332 373588
rect 563096 372880 563332 373116
rect 563096 372408 563332 372644
rect 563096 371936 563332 372172
rect 563096 371464 563332 371700
rect 563568 377128 563804 377364
rect 563568 376656 563804 376892
rect 563568 376184 563804 376420
rect 563568 375712 563804 375948
rect 563568 375240 563804 375476
rect 563568 374768 563804 375004
rect 563568 374296 563804 374532
rect 563568 373824 563804 374060
rect 563568 373352 563804 373588
rect 563568 372880 563804 373116
rect 563568 372408 563804 372644
rect 563568 371936 563804 372172
rect 563568 371464 563804 371700
rect 564040 377128 564276 377364
rect 564040 376656 564276 376892
rect 564040 376184 564276 376420
rect 564040 375712 564276 375948
rect 564040 375240 564276 375476
rect 564040 374768 564276 375004
rect 564040 374296 564276 374532
rect 564040 373824 564276 374060
rect 564040 373352 564276 373588
rect 564040 372880 564276 373116
rect 564040 372408 564276 372644
rect 564040 371936 564276 372172
rect 564040 371464 564276 371700
rect 564512 377128 564748 377364
rect 564512 376656 564748 376892
rect 564512 376184 564748 376420
rect 564512 375712 564748 375948
rect 564512 375240 564748 375476
rect 564512 374768 564748 375004
rect 564512 374296 564748 374532
rect 564512 373824 564748 374060
rect 564512 373352 564748 373588
rect 564512 372880 564748 373116
rect 564512 372408 564748 372644
rect 564512 371936 564748 372172
rect 564512 371464 564748 371700
rect 564984 377128 565220 377364
rect 564984 376656 565220 376892
rect 564984 376184 565220 376420
rect 564984 375712 565220 375948
rect 564984 375240 565220 375476
rect 564984 374768 565220 375004
rect 564984 374296 565220 374532
rect 564984 373824 565220 374060
rect 564984 373352 565220 373588
rect 564984 372880 565220 373116
rect 564984 372408 565220 372644
rect 564984 371936 565220 372172
rect 564984 371464 565220 371700
rect 565456 377128 565692 377364
rect 565456 376656 565692 376892
rect 565456 376184 565692 376420
rect 565456 375712 565692 375948
rect 565456 375240 565692 375476
rect 565456 374768 565692 375004
rect 565456 374296 565692 374532
rect 565456 373824 565692 374060
rect 565456 373352 565692 373588
rect 565456 372880 565692 373116
rect 565456 372408 565692 372644
rect 565456 371936 565692 372172
rect 565456 371464 565692 371700
rect 565928 377128 566164 377364
rect 565928 376656 566164 376892
rect 565928 376184 566164 376420
rect 565928 375712 566164 375948
rect 565928 375240 566164 375476
rect 565928 374768 566164 375004
rect 565928 374296 566164 374532
rect 565928 373824 566164 374060
rect 565928 373352 566164 373588
rect 565928 372880 566164 373116
rect 565928 372408 566164 372644
rect 565928 371936 566164 372172
rect 565928 371464 566164 371700
rect 566400 377128 566636 377364
rect 566400 376656 566636 376892
rect 566400 376184 566636 376420
rect 566400 375712 566636 375948
rect 566400 375240 566636 375476
rect 566400 374768 566636 375004
rect 566400 374296 566636 374532
rect 566400 373824 566636 374060
rect 566400 373352 566636 373588
rect 566400 372880 566636 373116
rect 566400 372408 566636 372644
rect 566400 371936 566636 372172
rect 566400 371464 566636 371700
rect 566872 377128 567108 377364
rect 566872 376656 567108 376892
rect 566872 376184 567108 376420
rect 566872 375712 567108 375948
rect 566872 375240 567108 375476
rect 566872 374768 567108 375004
rect 566872 374296 567108 374532
rect 566872 373824 567108 374060
rect 566872 373352 567108 373588
rect 566872 372880 567108 373116
rect 566872 372408 567108 372644
rect 566872 371936 567108 372172
rect 566872 371464 567108 371700
<< metal5 >>
rect 572560 697380 577480 697420
rect 572560 697144 577492 697380
rect 572560 696908 572772 697144
rect 573008 696908 573244 697144
rect 573480 696908 573716 697144
rect 573952 696908 574188 697144
rect 574424 696908 574660 697144
rect 574896 696908 575132 697144
rect 575368 696908 575604 697144
rect 575840 696908 576076 697144
rect 576312 696908 576548 697144
rect 576784 696908 577020 697144
rect 577256 696908 577492 697144
rect 572560 696672 577492 696908
rect 572560 696436 572772 696672
rect 573008 696436 573244 696672
rect 573480 696436 573716 696672
rect 573952 696436 574188 696672
rect 574424 696436 574660 696672
rect 574896 696436 575132 696672
rect 575368 696436 575604 696672
rect 575840 696436 576076 696672
rect 576312 696436 576548 696672
rect 576784 696436 577020 696672
rect 577256 696436 577492 696672
rect 572560 696200 577492 696436
rect 572560 695964 572772 696200
rect 573008 695964 573244 696200
rect 573480 695964 573716 696200
rect 573952 695964 574188 696200
rect 574424 695964 574660 696200
rect 574896 695964 575132 696200
rect 575368 695964 575604 696200
rect 575840 695964 576076 696200
rect 576312 695964 576548 696200
rect 576784 695964 577020 696200
rect 577256 695964 577492 696200
rect 572560 695728 577492 695964
rect 572560 695492 572772 695728
rect 573008 695492 573244 695728
rect 573480 695492 573716 695728
rect 573952 695492 574188 695728
rect 574424 695492 574660 695728
rect 574896 695492 575132 695728
rect 575368 695492 575604 695728
rect 575840 695492 576076 695728
rect 576312 695492 576548 695728
rect 576784 695492 577020 695728
rect 577256 695492 577492 695728
rect 572560 695256 577492 695492
rect 572560 695020 572772 695256
rect 573008 695020 573244 695256
rect 573480 695020 573716 695256
rect 573952 695020 574188 695256
rect 574424 695020 574660 695256
rect 574896 695020 575132 695256
rect 575368 695020 575604 695256
rect 575840 695020 576076 695256
rect 576312 695020 576548 695256
rect 576784 695020 577020 695256
rect 577256 695020 577492 695256
rect 572560 694784 577492 695020
rect 572560 694548 572772 694784
rect 573008 694548 573244 694784
rect 573480 694548 573716 694784
rect 573952 694548 574188 694784
rect 574424 694548 574660 694784
rect 574896 694548 575132 694784
rect 575368 694548 575604 694784
rect 575840 694548 576076 694784
rect 576312 694548 576548 694784
rect 576784 694548 577020 694784
rect 577256 694548 577492 694784
rect 572560 694312 577492 694548
rect 572560 694076 572772 694312
rect 573008 694076 573244 694312
rect 573480 694076 573716 694312
rect 573952 694076 574188 694312
rect 574424 694076 574660 694312
rect 574896 694076 575132 694312
rect 575368 694076 575604 694312
rect 575840 694076 576076 694312
rect 576312 694076 576548 694312
rect 576784 694076 577020 694312
rect 577256 694076 577492 694312
rect 572560 693840 577492 694076
rect 572560 693604 572772 693840
rect 573008 693604 573244 693840
rect 573480 693604 573716 693840
rect 573952 693604 574188 693840
rect 574424 693604 574660 693840
rect 574896 693604 575132 693840
rect 575368 693604 575604 693840
rect 575840 693604 576076 693840
rect 576312 693604 576548 693840
rect 576784 693604 577020 693840
rect 577256 693604 577492 693840
rect 572560 693368 577492 693604
rect 572560 693132 572772 693368
rect 573008 693132 573244 693368
rect 573480 693132 573716 693368
rect 573952 693132 574188 693368
rect 574424 693132 574660 693368
rect 574896 693132 575132 693368
rect 575368 693132 575604 693368
rect 575840 693132 576076 693368
rect 576312 693132 576548 693368
rect 576784 693132 577020 693368
rect 577256 693132 577492 693368
rect 572560 692896 577492 693132
rect 572560 692660 572772 692896
rect 573008 692660 573244 692896
rect 573480 692660 573716 692896
rect 573952 692660 574188 692896
rect 574424 692660 574660 692896
rect 574896 692660 575132 692896
rect 575368 692660 575604 692896
rect 575840 692660 576076 692896
rect 576312 692660 576548 692896
rect 576784 692660 577020 692896
rect 577256 692660 577492 692896
rect 562456 644584 567424 654608
rect 562456 639784 562480 644584
rect 567400 639784 567424 644584
rect 562456 634584 567424 639784
rect 562456 629784 562480 634584
rect 567400 629784 567424 634584
rect 562456 522504 567424 629784
rect 562456 522268 562624 522504
rect 562860 522268 563096 522504
rect 563332 522268 563568 522504
rect 563804 522268 564040 522504
rect 564276 522268 564512 522504
rect 564748 522268 564984 522504
rect 565220 522268 565456 522504
rect 565692 522268 565928 522504
rect 566164 522268 566400 522504
rect 566636 522268 566872 522504
rect 567108 522268 567424 522504
rect 562456 522032 567424 522268
rect 562456 521796 562624 522032
rect 562860 521796 563096 522032
rect 563332 521796 563568 522032
rect 563804 521796 564040 522032
rect 564276 521796 564512 522032
rect 564748 521796 564984 522032
rect 565220 521796 565456 522032
rect 565692 521796 565928 522032
rect 566164 521796 566400 522032
rect 566636 521796 566872 522032
rect 567108 521796 567424 522032
rect 562456 521560 567424 521796
rect 562456 521324 562624 521560
rect 562860 521324 563096 521560
rect 563332 521324 563568 521560
rect 563804 521324 564040 521560
rect 564276 521324 564512 521560
rect 564748 521324 564984 521560
rect 565220 521324 565456 521560
rect 565692 521324 565928 521560
rect 566164 521324 566400 521560
rect 566636 521324 566872 521560
rect 567108 521324 567424 521560
rect 562456 521088 567424 521324
rect 562456 520852 562624 521088
rect 562860 520852 563096 521088
rect 563332 520852 563568 521088
rect 563804 520852 564040 521088
rect 564276 520852 564512 521088
rect 564748 520852 564984 521088
rect 565220 520852 565456 521088
rect 565692 520852 565928 521088
rect 566164 520852 566400 521088
rect 566636 520852 566872 521088
rect 567108 520852 567424 521088
rect 562456 520616 567424 520852
rect 562456 520380 562624 520616
rect 562860 520380 563096 520616
rect 563332 520380 563568 520616
rect 563804 520380 564040 520616
rect 564276 520380 564512 520616
rect 564748 520380 564984 520616
rect 565220 520380 565456 520616
rect 565692 520380 565928 520616
rect 566164 520380 566400 520616
rect 566636 520380 566872 520616
rect 567108 520380 567424 520616
rect 562456 520144 567424 520380
rect 562456 519908 562624 520144
rect 562860 519908 563096 520144
rect 563332 519908 563568 520144
rect 563804 519908 564040 520144
rect 564276 519908 564512 520144
rect 564748 519908 564984 520144
rect 565220 519908 565456 520144
rect 565692 519908 565928 520144
rect 566164 519908 566400 520144
rect 566636 519908 566872 520144
rect 567108 519908 567424 520144
rect 562456 519672 567424 519908
rect 562456 519436 562624 519672
rect 562860 519436 563096 519672
rect 563332 519436 563568 519672
rect 563804 519436 564040 519672
rect 564276 519436 564512 519672
rect 564748 519436 564984 519672
rect 565220 519436 565456 519672
rect 565692 519436 565928 519672
rect 566164 519436 566400 519672
rect 566636 519436 566872 519672
rect 567108 519436 567424 519672
rect 562456 519200 567424 519436
rect 562456 518964 562624 519200
rect 562860 518964 563096 519200
rect 563332 518964 563568 519200
rect 563804 518964 564040 519200
rect 564276 518964 564512 519200
rect 564748 518964 564984 519200
rect 565220 518964 565456 519200
rect 565692 518964 565928 519200
rect 566164 518964 566400 519200
rect 566636 518964 566872 519200
rect 567108 518964 567424 519200
rect 562456 518728 567424 518964
rect 562456 518492 562624 518728
rect 562860 518492 563096 518728
rect 563332 518492 563568 518728
rect 563804 518492 564040 518728
rect 564276 518492 564512 518728
rect 564748 518492 564984 518728
rect 565220 518492 565456 518728
rect 565692 518492 565928 518728
rect 566164 518492 566400 518728
rect 566636 518492 566872 518728
rect 567108 518492 567424 518728
rect 562456 518256 567424 518492
rect 562456 518020 562624 518256
rect 562860 518020 563096 518256
rect 563332 518020 563568 518256
rect 563804 518020 564040 518256
rect 564276 518020 564512 518256
rect 564748 518020 564984 518256
rect 565220 518020 565456 518256
rect 565692 518020 565928 518256
rect 566164 518020 566400 518256
rect 566636 518020 566872 518256
rect 567108 518020 567424 518256
rect 562456 517784 567424 518020
rect 562456 517548 562624 517784
rect 562860 517548 563096 517784
rect 563332 517548 563568 517784
rect 563804 517548 564040 517784
rect 564276 517548 564512 517784
rect 564748 517548 564984 517784
rect 565220 517548 565456 517784
rect 565692 517548 565928 517784
rect 566164 517548 566400 517784
rect 566636 517548 566872 517784
rect 567108 517548 567424 517784
rect 562456 517312 567424 517548
rect 562456 517076 562624 517312
rect 562860 517076 563096 517312
rect 563332 517076 563568 517312
rect 563804 517076 564040 517312
rect 564276 517076 564512 517312
rect 564748 517076 564984 517312
rect 565220 517076 565456 517312
rect 565692 517076 565928 517312
rect 566164 517076 566400 517312
rect 566636 517076 566872 517312
rect 567108 517076 567424 517312
rect 562456 516840 567424 517076
rect 562456 516604 562624 516840
rect 562860 516604 563096 516840
rect 563332 516604 563568 516840
rect 563804 516604 564040 516840
rect 564276 516604 564512 516840
rect 564748 516604 564984 516840
rect 565220 516604 565456 516840
rect 565692 516604 565928 516840
rect 566164 516604 566400 516840
rect 566636 516604 566872 516840
rect 567108 516604 567424 516840
rect 562456 495782 567424 516604
rect 562456 495546 562624 495782
rect 562860 495546 563096 495782
rect 563332 495546 563568 495782
rect 563804 495546 564040 495782
rect 564276 495546 564512 495782
rect 564748 495546 564984 495782
rect 565220 495546 565456 495782
rect 565692 495546 565928 495782
rect 566164 495546 566400 495782
rect 566636 495546 566872 495782
rect 567108 495546 567424 495782
rect 562456 455480 567424 495546
rect 562456 455244 562624 455480
rect 562860 455244 563096 455480
rect 563332 455244 563568 455480
rect 563804 455244 564040 455480
rect 564276 455244 564512 455480
rect 564748 455244 564984 455480
rect 565220 455244 565456 455480
rect 565692 455244 565928 455480
rect 566164 455244 566400 455480
rect 566636 455244 566872 455480
rect 567108 455244 567424 455480
rect 562456 377364 567424 455244
rect 562456 377128 562624 377364
rect 562860 377128 563096 377364
rect 563332 377128 563568 377364
rect 563804 377128 564040 377364
rect 564276 377128 564512 377364
rect 564748 377128 564984 377364
rect 565220 377128 565456 377364
rect 565692 377128 565928 377364
rect 566164 377128 566400 377364
rect 566636 377128 566872 377364
rect 567108 377128 567424 377364
rect 562456 376892 567424 377128
rect 562456 376656 562624 376892
rect 562860 376656 563096 376892
rect 563332 376656 563568 376892
rect 563804 376656 564040 376892
rect 564276 376656 564512 376892
rect 564748 376656 564984 376892
rect 565220 376656 565456 376892
rect 565692 376656 565928 376892
rect 566164 376656 566400 376892
rect 566636 376656 566872 376892
rect 567108 376656 567424 376892
rect 562456 376420 567424 376656
rect 562456 376184 562624 376420
rect 562860 376184 563096 376420
rect 563332 376184 563568 376420
rect 563804 376184 564040 376420
rect 564276 376184 564512 376420
rect 564748 376184 564984 376420
rect 565220 376184 565456 376420
rect 565692 376184 565928 376420
rect 566164 376184 566400 376420
rect 566636 376184 566872 376420
rect 567108 376184 567424 376420
rect 562456 375948 567424 376184
rect 562456 375712 562624 375948
rect 562860 375712 563096 375948
rect 563332 375712 563568 375948
rect 563804 375712 564040 375948
rect 564276 375712 564512 375948
rect 564748 375712 564984 375948
rect 565220 375712 565456 375948
rect 565692 375712 565928 375948
rect 566164 375712 566400 375948
rect 566636 375712 566872 375948
rect 567108 375712 567424 375948
rect 562456 375476 567424 375712
rect 562456 375240 562624 375476
rect 562860 375240 563096 375476
rect 563332 375240 563568 375476
rect 563804 375240 564040 375476
rect 564276 375240 564512 375476
rect 564748 375240 564984 375476
rect 565220 375240 565456 375476
rect 565692 375240 565928 375476
rect 566164 375240 566400 375476
rect 566636 375240 566872 375476
rect 567108 375240 567424 375476
rect 562456 375004 567424 375240
rect 562456 374768 562624 375004
rect 562860 374768 563096 375004
rect 563332 374768 563568 375004
rect 563804 374768 564040 375004
rect 564276 374768 564512 375004
rect 564748 374768 564984 375004
rect 565220 374768 565456 375004
rect 565692 374768 565928 375004
rect 566164 374768 566400 375004
rect 566636 374768 566872 375004
rect 567108 374768 567424 375004
rect 562456 374532 567424 374768
rect 562456 374296 562624 374532
rect 562860 374296 563096 374532
rect 563332 374296 563568 374532
rect 563804 374296 564040 374532
rect 564276 374296 564512 374532
rect 564748 374296 564984 374532
rect 565220 374296 565456 374532
rect 565692 374296 565928 374532
rect 566164 374296 566400 374532
rect 566636 374296 566872 374532
rect 567108 374296 567424 374532
rect 562456 374060 567424 374296
rect 562456 373824 562624 374060
rect 562860 373824 563096 374060
rect 563332 373824 563568 374060
rect 563804 373824 564040 374060
rect 564276 373824 564512 374060
rect 564748 373824 564984 374060
rect 565220 373824 565456 374060
rect 565692 373824 565928 374060
rect 566164 373824 566400 374060
rect 566636 373824 566872 374060
rect 567108 373824 567424 374060
rect 562456 373588 567424 373824
rect 562456 373352 562624 373588
rect 562860 373352 563096 373588
rect 563332 373352 563568 373588
rect 563804 373352 564040 373588
rect 564276 373352 564512 373588
rect 564748 373352 564984 373588
rect 565220 373352 565456 373588
rect 565692 373352 565928 373588
rect 566164 373352 566400 373588
rect 566636 373352 566872 373588
rect 567108 373352 567424 373588
rect 562456 373116 567424 373352
rect 562456 372880 562624 373116
rect 562860 372880 563096 373116
rect 563332 372880 563568 373116
rect 563804 372880 564040 373116
rect 564276 372880 564512 373116
rect 564748 372880 564984 373116
rect 565220 372880 565456 373116
rect 565692 372880 565928 373116
rect 566164 372880 566400 373116
rect 566636 372880 566872 373116
rect 567108 372880 567424 373116
rect 562456 372644 567424 372880
rect 562456 372408 562624 372644
rect 562860 372408 563096 372644
rect 563332 372408 563568 372644
rect 563804 372408 564040 372644
rect 564276 372408 564512 372644
rect 564748 372408 564984 372644
rect 565220 372408 565456 372644
rect 565692 372408 565928 372644
rect 566164 372408 566400 372644
rect 566636 372408 566872 372644
rect 567108 372408 567424 372644
rect 562456 372172 567424 372408
rect 562456 371936 562624 372172
rect 562860 371936 563096 372172
rect 563332 371936 563568 372172
rect 563804 371936 564040 372172
rect 564276 371936 564512 372172
rect 564748 371936 564984 372172
rect 565220 371936 565456 372172
rect 565692 371936 565928 372172
rect 566164 371936 566400 372172
rect 566636 371936 566872 372172
rect 567108 371936 567424 372172
rect 562456 371700 567424 371936
rect 562456 371464 562624 371700
rect 562860 371464 563096 371700
rect 563332 371464 563568 371700
rect 563804 371464 564040 371700
rect 564276 371464 564512 371700
rect 564748 371464 564984 371700
rect 565220 371464 565456 371700
rect 565692 371464 565928 371700
rect 566164 371464 566400 371700
rect 566636 371464 566872 371700
rect 567108 371464 567424 371700
rect 562456 303322 567424 371464
rect 572560 495782 577480 692660
rect 572560 495546 572784 495782
rect 573020 495546 573256 495782
rect 573492 495546 573728 495782
rect 573964 495546 574200 495782
rect 574436 495546 574672 495782
rect 574908 495546 575144 495782
rect 575380 495546 575616 495782
rect 575852 495546 576088 495782
rect 576324 495546 576560 495782
rect 576796 495546 577032 495782
rect 577268 495546 577480 495782
rect 572560 484272 577480 495546
rect 572560 484036 577492 484272
rect 572560 483800 572772 484036
rect 573008 483800 573244 484036
rect 573480 483800 573716 484036
rect 573952 483800 574188 484036
rect 574424 483800 574660 484036
rect 574896 483800 575132 484036
rect 575368 483800 575604 484036
rect 575840 483800 576076 484036
rect 576312 483800 576548 484036
rect 576784 483800 577020 484036
rect 577256 483800 577492 484036
rect 572560 483564 577492 483800
rect 572560 483328 572772 483564
rect 573008 483328 573244 483564
rect 573480 483328 573716 483564
rect 573952 483328 574188 483564
rect 574424 483328 574660 483564
rect 574896 483328 575132 483564
rect 575368 483328 575604 483564
rect 575840 483328 576076 483564
rect 576312 483328 576548 483564
rect 576784 483328 577020 483564
rect 577256 483328 577492 483564
rect 572560 483092 577492 483328
rect 572560 482856 572772 483092
rect 573008 482856 573244 483092
rect 573480 482856 573716 483092
rect 573952 482856 574188 483092
rect 574424 482856 574660 483092
rect 574896 482856 575132 483092
rect 575368 482856 575604 483092
rect 575840 482856 576076 483092
rect 576312 482856 576548 483092
rect 576784 482856 577020 483092
rect 577256 482856 577492 483092
rect 572560 482620 577492 482856
rect 572560 482384 572772 482620
rect 573008 482384 573244 482620
rect 573480 482384 573716 482620
rect 573952 482384 574188 482620
rect 574424 482384 574660 482620
rect 574896 482384 575132 482620
rect 575368 482384 575604 482620
rect 575840 482384 576076 482620
rect 576312 482384 576548 482620
rect 576784 482384 577020 482620
rect 577256 482384 577492 482620
rect 572560 482148 577492 482384
rect 572560 481912 572772 482148
rect 573008 481912 573244 482148
rect 573480 481912 573716 482148
rect 573952 481912 574188 482148
rect 574424 481912 574660 482148
rect 574896 481912 575132 482148
rect 575368 481912 575604 482148
rect 575840 481912 576076 482148
rect 576312 481912 576548 482148
rect 576784 481912 577020 482148
rect 577256 481912 577492 482148
rect 572560 481676 577492 481912
rect 572560 481440 572772 481676
rect 573008 481440 573244 481676
rect 573480 481440 573716 481676
rect 573952 481440 574188 481676
rect 574424 481440 574660 481676
rect 574896 481440 575132 481676
rect 575368 481440 575604 481676
rect 575840 481440 576076 481676
rect 576312 481440 576548 481676
rect 576784 481440 577020 481676
rect 577256 481440 577492 481676
rect 572560 481204 577492 481440
rect 572560 480968 572772 481204
rect 573008 480968 573244 481204
rect 573480 480968 573716 481204
rect 573952 480968 574188 481204
rect 574424 480968 574660 481204
rect 574896 480968 575132 481204
rect 575368 480968 575604 481204
rect 575840 480968 576076 481204
rect 576312 480968 576548 481204
rect 576784 480968 577020 481204
rect 577256 480968 577492 481204
rect 572560 480732 577492 480968
rect 572560 480496 572772 480732
rect 573008 480496 573244 480732
rect 573480 480496 573716 480732
rect 573952 480496 574188 480732
rect 574424 480496 574660 480732
rect 574896 480496 575132 480732
rect 575368 480496 575604 480732
rect 575840 480496 576076 480732
rect 576312 480496 576548 480732
rect 576784 480496 577020 480732
rect 577256 480496 577492 480732
rect 572560 480260 577492 480496
rect 572560 480024 572772 480260
rect 573008 480024 573244 480260
rect 573480 480024 573716 480260
rect 573952 480024 574188 480260
rect 574424 480024 574660 480260
rect 574896 480024 575132 480260
rect 575368 480024 575604 480260
rect 575840 480024 576076 480260
rect 576312 480024 576548 480260
rect 576784 480024 577020 480260
rect 577256 480024 577492 480260
rect 572560 479788 577492 480024
rect 572560 479552 572772 479788
rect 573008 479552 573244 479788
rect 573480 479552 573716 479788
rect 573952 479552 574188 479788
rect 574424 479552 574660 479788
rect 574896 479552 575132 479788
rect 575368 479552 575604 479788
rect 575840 479552 576076 479788
rect 576312 479552 576548 479788
rect 576784 479552 577020 479788
rect 577256 479552 577492 479788
rect 572560 479316 577492 479552
rect 572560 479080 572772 479316
rect 573008 479080 573244 479316
rect 573480 479080 573716 479316
rect 573952 479080 574188 479316
rect 574424 479080 574660 479316
rect 574896 479080 575132 479316
rect 575368 479080 575604 479316
rect 575840 479080 576076 479316
rect 576312 479080 576548 479316
rect 576784 479080 577020 479316
rect 577256 479080 577492 479316
rect 572560 478844 577492 479080
rect 572560 478608 572772 478844
rect 573008 478608 573244 478844
rect 573480 478608 573716 478844
rect 573952 478608 574188 478844
rect 574424 478608 574660 478844
rect 574896 478608 575132 478844
rect 575368 478608 575604 478844
rect 575840 478608 576076 478844
rect 576312 478608 576548 478844
rect 576784 478608 577020 478844
rect 577256 478608 577492 478844
rect 572560 478372 577492 478608
rect 572560 478136 572772 478372
rect 573008 478136 573244 478372
rect 573480 478136 573716 478372
rect 573952 478136 574188 478372
rect 574424 478136 574660 478372
rect 574896 478136 575132 478372
rect 575368 478136 575604 478372
rect 575840 478136 576076 478372
rect 576312 478136 576548 478372
rect 576784 478136 577020 478372
rect 577256 478136 577492 478372
rect 572560 477900 577492 478136
rect 572560 477664 572772 477900
rect 573008 477664 573244 477900
rect 573480 477664 573716 477900
rect 573952 477664 574188 477900
rect 574424 477664 574660 477900
rect 574896 477664 575132 477900
rect 575368 477664 575604 477900
rect 575840 477664 576076 477900
rect 576312 477664 576548 477900
rect 576784 477664 577020 477900
rect 577256 477664 577492 477900
rect 572560 455480 577480 477664
rect 572560 455244 572784 455480
rect 573020 455244 573256 455480
rect 573492 455244 573728 455480
rect 573964 455244 574200 455480
rect 574436 455244 574672 455480
rect 574908 455244 575144 455480
rect 575380 455244 575616 455480
rect 575852 455244 576088 455480
rect 576324 455244 576560 455480
rect 576796 455244 577032 455480
rect 577268 455244 577480 455480
rect 572560 426924 577480 455244
rect 572560 426688 577492 426924
rect 572560 426452 572772 426688
rect 573008 426452 573244 426688
rect 573480 426452 573716 426688
rect 573952 426452 574188 426688
rect 574424 426452 574660 426688
rect 574896 426452 575132 426688
rect 575368 426452 575604 426688
rect 575840 426452 576076 426688
rect 576312 426452 576548 426688
rect 576784 426452 577020 426688
rect 577256 426452 577492 426688
rect 572560 426216 577492 426452
rect 572560 425980 572772 426216
rect 573008 425980 573244 426216
rect 573480 425980 573716 426216
rect 573952 425980 574188 426216
rect 574424 425980 574660 426216
rect 574896 425980 575132 426216
rect 575368 425980 575604 426216
rect 575840 425980 576076 426216
rect 576312 425980 576548 426216
rect 576784 425980 577020 426216
rect 577256 425980 577492 426216
rect 572560 425744 577492 425980
rect 572560 425508 572772 425744
rect 573008 425508 573244 425744
rect 573480 425508 573716 425744
rect 573952 425508 574188 425744
rect 574424 425508 574660 425744
rect 574896 425508 575132 425744
rect 575368 425508 575604 425744
rect 575840 425508 576076 425744
rect 576312 425508 576548 425744
rect 576784 425508 577020 425744
rect 577256 425508 577492 425744
rect 572560 425272 577492 425508
rect 572560 425036 572772 425272
rect 573008 425036 573244 425272
rect 573480 425036 573716 425272
rect 573952 425036 574188 425272
rect 574424 425036 574660 425272
rect 574896 425036 575132 425272
rect 575368 425036 575604 425272
rect 575840 425036 576076 425272
rect 576312 425036 576548 425272
rect 576784 425036 577020 425272
rect 577256 425036 577492 425272
rect 572560 424800 577492 425036
rect 572560 424564 572772 424800
rect 573008 424564 573244 424800
rect 573480 424564 573716 424800
rect 573952 424564 574188 424800
rect 574424 424564 574660 424800
rect 574896 424564 575132 424800
rect 575368 424564 575604 424800
rect 575840 424564 576076 424800
rect 576312 424564 576548 424800
rect 576784 424564 577020 424800
rect 577256 424564 577492 424800
rect 572560 424328 577492 424564
rect 572560 424092 572772 424328
rect 573008 424092 573244 424328
rect 573480 424092 573716 424328
rect 573952 424092 574188 424328
rect 574424 424092 574660 424328
rect 574896 424092 575132 424328
rect 575368 424092 575604 424328
rect 575840 424092 576076 424328
rect 576312 424092 576548 424328
rect 576784 424092 577020 424328
rect 577256 424092 577492 424328
rect 572560 423856 577492 424092
rect 572560 423620 572772 423856
rect 573008 423620 573244 423856
rect 573480 423620 573716 423856
rect 573952 423620 574188 423856
rect 574424 423620 574660 423856
rect 574896 423620 575132 423856
rect 575368 423620 575604 423856
rect 575840 423620 576076 423856
rect 576312 423620 576548 423856
rect 576784 423620 577020 423856
rect 577256 423620 577492 423856
rect 572560 423384 577492 423620
rect 572560 423148 572772 423384
rect 573008 423148 573244 423384
rect 573480 423148 573716 423384
rect 573952 423148 574188 423384
rect 574424 423148 574660 423384
rect 574896 423148 575132 423384
rect 575368 423148 575604 423384
rect 575840 423148 576076 423384
rect 576312 423148 576548 423384
rect 576784 423148 577020 423384
rect 577256 423148 577492 423384
rect 572560 422912 577492 423148
rect 572560 422676 572772 422912
rect 573008 422676 573244 422912
rect 573480 422676 573716 422912
rect 573952 422676 574188 422912
rect 574424 422676 574660 422912
rect 574896 422676 575132 422912
rect 575368 422676 575604 422912
rect 575840 422676 576076 422912
rect 576312 422676 576548 422912
rect 576784 422676 577020 422912
rect 577256 422676 577492 422912
rect 572560 422440 577492 422676
rect 572560 422204 572772 422440
rect 573008 422204 573244 422440
rect 573480 422204 573716 422440
rect 573952 422204 574188 422440
rect 574424 422204 574660 422440
rect 574896 422204 575132 422440
rect 575368 422204 575604 422440
rect 575840 422204 576076 422440
rect 576312 422204 576548 422440
rect 576784 422204 577020 422440
rect 577256 422204 577492 422440
rect 572560 421968 577492 422204
rect 572560 421732 572772 421968
rect 573008 421732 573244 421968
rect 573480 421732 573716 421968
rect 573952 421732 574188 421968
rect 574424 421732 574660 421968
rect 574896 421732 575132 421968
rect 575368 421732 575604 421968
rect 575840 421732 576076 421968
rect 576312 421732 576548 421968
rect 576784 421732 577020 421968
rect 577256 421732 577492 421968
rect 572560 421496 577492 421732
rect 572560 421260 572772 421496
rect 573008 421260 573244 421496
rect 573480 421260 573716 421496
rect 573952 421260 574188 421496
rect 574424 421260 574660 421496
rect 574896 421260 575132 421496
rect 575368 421260 575604 421496
rect 575840 421260 576076 421496
rect 576312 421260 576548 421496
rect 576784 421260 577020 421496
rect 577256 421260 577492 421496
rect 572560 421024 577492 421260
rect 572560 420788 572772 421024
rect 573008 420788 573244 421024
rect 573480 420788 573716 421024
rect 573952 420788 574188 421024
rect 574424 420788 574660 421024
rect 574896 420788 575132 421024
rect 575368 420788 575604 421024
rect 575840 420788 576076 421024
rect 576312 420788 576548 421024
rect 576784 420788 577020 421024
rect 577256 420788 577492 421024
rect 572560 420552 577492 420788
rect 572560 420316 572772 420552
rect 573008 420316 573244 420552
rect 573480 420316 573716 420552
rect 573952 420316 574188 420552
rect 574424 420316 574660 420552
rect 574896 420316 575132 420552
rect 575368 420316 575604 420552
rect 575840 420316 576076 420552
rect 576312 420316 576548 420552
rect 576784 420316 577020 420552
rect 577256 420316 577492 420552
rect 572560 312500 577480 420316
<< comment >>
rect -100 704000 584100 704100
rect -100 0 0 704000
rect 584000 0 584100 704000
rect -100 -100 584100 0
use sky130_fd_pr__nfet_01v8_lvt_ZQXVKQ  sky130_fd_pr__nfet_01v8_lvt_ZQXVKQ_1
timestamp 1622316573
transform 1 0 575027 0 -1 494905
box -2747 -679 2747 679
use sky130_fd_pr__pfet_01v8_lvt_V33E7D  sky130_fd_pr__pfet_01v8_lvt_V33E7D_1
timestamp 1622314978
transform -1 0 564867 0 -1 494866
box -2747 -684 2747 684
use bandgaptop_flat_io  bandgaptop_flat_io_0
timestamp 1622225665
transform 0 1 -126262 -1 0 913200
box 422960 603262 502000 669400
use sky130_fd_pr__pfet_01v8_lvt_V33E7D  sky130_fd_pr__pfet_01v8_lvt_V33E7D_0
timestamp 1622314978
transform -1 0 564867 0 -1 454564
box -2747 -684 2747 684
use sky130_fd_pr__nfet_01v8_lvt_ZQXVKQ  sky130_fd_pr__nfet_01v8_lvt_ZQXVKQ_0
timestamp 1622316573
transform 1 0 575027 0 -1 454603
box -2747 -679 2747 679
<< labels >>
flabel metal3 s 583520 269230 584800 269342 0 FreeSans 1120 0 0 0 gpio_analog[0]
port 0 nsew signal bidirectional
flabel metal3 s -800 381864 480 381976 0 FreeSans 1120 0 0 0 gpio_analog[10]
port 1 nsew signal bidirectional
flabel metal3 s -800 338642 480 338754 0 FreeSans 1120 0 0 0 gpio_analog[11]
port 2 nsew signal bidirectional
flabel metal3 s -800 295420 480 295532 0 FreeSans 1120 0 0 0 gpio_analog[12]
port 3 nsew signal bidirectional
flabel metal3 s -800 252398 480 252510 0 FreeSans 1120 0 0 0 gpio_analog[13]
port 4 nsew signal bidirectional
flabel metal3 s -800 124776 480 124888 0 FreeSans 1120 0 0 0 gpio_analog[14]
port 5 nsew signal bidirectional
flabel metal3 s -800 81554 480 81666 0 FreeSans 1120 0 0 0 gpio_analog[15]
port 6 nsew signal bidirectional
flabel metal3 s -800 38332 480 38444 0 FreeSans 1120 0 0 0 gpio_analog[16]
port 7 nsew signal bidirectional
flabel metal3 s -800 16910 480 17022 0 FreeSans 1120 0 0 0 gpio_analog[17]
port 8 nsew signal bidirectional
flabel metal3 s 583520 313652 584800 313764 0 FreeSans 1120 0 0 0 gpio_analog[1]
port 9 nsew signal bidirectional
flabel metal3 s 583520 358874 584800 358986 0 FreeSans 1120 0 0 0 gpio_analog[2]
port 10 nsew signal bidirectional
flabel metal3 s 583520 405296 584800 405408 0 FreeSans 1120 0 0 0 gpio_analog[3]
port 11 nsew signal bidirectional
flabel metal3 s 583520 449718 584800 449830 0 FreeSans 1120 0 0 0 gpio_analog[4]
port 12 nsew signal bidirectional
flabel metal3 s 583520 494140 584800 494252 0 FreeSans 1120 0 0 0 gpio_analog[5]
port 13 nsew signal bidirectional
flabel metal3 s 583520 583562 584800 583674 0 FreeSans 1120 0 0 0 gpio_analog[6]
port 14 nsew signal bidirectional
flabel metal3 s -800 511530 480 511642 0 FreeSans 1120 0 0 0 gpio_analog[7]
port 15 nsew signal bidirectional
flabel metal3 s -800 468308 480 468420 0 FreeSans 1120 0 0 0 gpio_analog[8]
port 16 nsew signal bidirectional
flabel metal3 s -800 425086 480 425198 0 FreeSans 1120 0 0 0 gpio_analog[9]
port 17 nsew signal bidirectional
flabel metal3 s 583520 270412 584800 270524 0 FreeSans 1120 0 0 0 gpio_noesd[0]
port 18 nsew signal bidirectional
flabel metal3 s -800 380682 480 380794 0 FreeSans 1120 0 0 0 gpio_noesd[10]
port 19 nsew signal bidirectional
flabel metal3 s -800 337460 480 337572 0 FreeSans 1120 0 0 0 gpio_noesd[11]
port 20 nsew signal bidirectional
flabel metal3 s -800 294238 480 294350 0 FreeSans 1120 0 0 0 gpio_noesd[12]
port 21 nsew signal bidirectional
flabel metal3 s -800 251216 480 251328 0 FreeSans 1120 0 0 0 gpio_noesd[13]
port 22 nsew signal bidirectional
flabel metal3 s -800 123594 480 123706 0 FreeSans 1120 0 0 0 gpio_noesd[14]
port 23 nsew signal bidirectional
flabel metal3 s -800 80372 480 80484 0 FreeSans 1120 0 0 0 gpio_noesd[15]
port 24 nsew signal bidirectional
flabel metal3 s -800 37150 480 37262 0 FreeSans 1120 0 0 0 gpio_noesd[16]
port 25 nsew signal bidirectional
flabel metal3 s -800 15728 480 15840 0 FreeSans 1120 0 0 0 gpio_noesd[17]
port 26 nsew signal bidirectional
flabel metal3 s 583520 314834 584800 314946 0 FreeSans 1120 0 0 0 gpio_noesd[1]
port 27 nsew signal bidirectional
flabel metal3 s 583520 360056 584800 360168 0 FreeSans 1120 0 0 0 gpio_noesd[2]
port 28 nsew signal bidirectional
flabel metal3 s 583520 406478 584800 406590 0 FreeSans 1120 0 0 0 gpio_noesd[3]
port 29 nsew signal bidirectional
flabel metal3 s 583520 450900 584800 451012 0 FreeSans 1120 0 0 0 gpio_noesd[4]
port 30 nsew signal bidirectional
flabel metal3 s 583520 495322 584800 495434 0 FreeSans 1120 0 0 0 gpio_noesd[5]
port 31 nsew signal bidirectional
flabel metal3 s 583520 584744 584800 584856 0 FreeSans 1120 0 0 0 gpio_noesd[6]
port 32 nsew signal bidirectional
flabel metal3 s -800 510348 480 510460 0 FreeSans 1120 0 0 0 gpio_noesd[7]
port 33 nsew signal bidirectional
flabel metal3 s -800 467126 480 467238 0 FreeSans 1120 0 0 0 gpio_noesd[8]
port 34 nsew signal bidirectional
flabel metal3 s -800 423904 480 424016 0 FreeSans 1120 0 0 0 gpio_noesd[9]
port 35 nsew signal bidirectional
flabel metal3 s 582300 677984 584800 682984 0 FreeSans 1120 0 0 0 io_analog[0]
port 36 nsew signal bidirectional
flabel metal3 s 0 680242 1700 685242 0 FreeSans 1120 0 0 0 io_analog[10]
port 37 nsew signal bidirectional
flabel metal3 s 566594 702300 571594 704800 0 FreeSans 1920 180 0 0 io_analog[1]
port 38 nsew signal bidirectional
flabel metal3 s 465394 702300 470394 704800 0 FreeSans 1920 180 0 0 io_analog[2]
port 39 nsew signal bidirectional
flabel metal3 s 413394 702300 418394 704800 0 FreeSans 1920 180 0 0 io_analog[3]
port 40 nsew signal bidirectional
flabel metal3 s 329294 702300 334294 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 41 nsew signal bidirectional
flabel metal3 s 227594 702300 232594 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 42 nsew signal bidirectional
flabel metal3 s 175894 702300 180894 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 43 nsew signal bidirectional
flabel metal3 s 120194 702300 125194 704800 0 FreeSans 1920 180 0 0 io_analog[7]
port 44 nsew signal bidirectional
flabel metal3 s 68194 702300 73194 704800 0 FreeSans 1920 180 0 0 io_analog[8]
port 45 nsew signal bidirectional
flabel metal3 s 16194 702300 21194 704800 0 FreeSans 1920 180 0 0 io_analog[9]
port 46 nsew signal bidirectional
flabel metal3 s 318994 702300 323994 704800 0 FreeSans 1920 180 0 0 io_analog[4]
port 47 nsew signal bidirectional
flabel metal3 s 217294 702300 222294 704800 0 FreeSans 1920 180 0 0 io_analog[5]
port 48 nsew signal bidirectional
flabel metal3 s 165594 702300 170594 704800 0 FreeSans 1920 180 0 0 io_analog[6]
port 49 nsew signal bidirectional
flabel metal3 s 326794 702300 328994 704800 0 FreeSans 1920 180 0 0 io_clamp_high[0]
port 50 nsew signal bidirectional
flabel metal3 s 225094 702300 227294 704800 0 FreeSans 1920 180 0 0 io_clamp_high[1]
port 51 nsew signal bidirectional
flabel metal3 s 173394 702300 175594 704800 0 FreeSans 1920 180 0 0 io_clamp_high[2]
port 52 nsew signal bidirectional
flabel metal3 s 324294 702300 326494 704800 0 FreeSans 1920 180 0 0 io_clamp_low[0]
port 53 nsew signal bidirectional
flabel metal3 s 222594 702300 224794 704800 0 FreeSans 1920 180 0 0 io_clamp_low[1]
port 54 nsew signal bidirectional
flabel metal3 s 170894 702300 173094 704800 0 FreeSans 1920 180 0 0 io_clamp_low[2]
port 55 nsew signal bidirectional
flabel metal3 s 583520 2726 584800 2838 0 FreeSans 1120 0 0 0 io_in[0]
port 56 nsew signal input
flabel metal3 s 583520 408842 584800 408954 0 FreeSans 1120 0 0 0 io_in[10]
port 57 nsew signal input
flabel metal3 s 583520 453264 584800 453376 0 FreeSans 1120 0 0 0 io_in[11]
port 58 nsew signal input
flabel metal3 s 583520 497686 584800 497798 0 FreeSans 1120 0 0 0 io_in[12]
port 59 nsew signal input
flabel metal3 s 583520 587108 584800 587220 0 FreeSans 1120 0 0 0 io_in[13]
port 60 nsew signal input
flabel metal3 s -800 507984 480 508096 0 FreeSans 1120 0 0 0 io_in[14]
port 61 nsew signal input
flabel metal3 s -800 464762 480 464874 0 FreeSans 1120 0 0 0 io_in[15]
port 62 nsew signal input
flabel metal3 s -800 421540 480 421652 0 FreeSans 1120 0 0 0 io_in[16]
port 63 nsew signal input
flabel metal3 s -800 378318 480 378430 0 FreeSans 1120 0 0 0 io_in[17]
port 64 nsew signal input
flabel metal3 s -800 335096 480 335208 0 FreeSans 1120 0 0 0 io_in[18]
port 65 nsew signal input
flabel metal3 s -800 291874 480 291986 0 FreeSans 1120 0 0 0 io_in[19]
port 66 nsew signal input
flabel metal3 s 583520 7454 584800 7566 0 FreeSans 1120 0 0 0 io_in[1]
port 67 nsew signal input
flabel metal3 s -800 248852 480 248964 0 FreeSans 1120 0 0 0 io_in[20]
port 68 nsew signal input
flabel metal3 s -800 121230 480 121342 0 FreeSans 1120 0 0 0 io_in[21]
port 69 nsew signal input
flabel metal3 s -800 78008 480 78120 0 FreeSans 1120 0 0 0 io_in[22]
port 70 nsew signal input
flabel metal3 s -800 34786 480 34898 0 FreeSans 1120 0 0 0 io_in[23]
port 71 nsew signal input
flabel metal3 s -800 13364 480 13476 0 FreeSans 1120 0 0 0 io_in[24]
port 72 nsew signal input
flabel metal3 s -800 8636 480 8748 0 FreeSans 1120 0 0 0 io_in[25]
port 73 nsew signal input
flabel metal3 s -800 3908 480 4020 0 FreeSans 1120 0 0 0 io_in[26]
port 74 nsew signal input
flabel metal3 s 583520 12182 584800 12294 0 FreeSans 1120 0 0 0 io_in[2]
port 75 nsew signal input
flabel metal3 s 583520 16910 584800 17022 0 FreeSans 1120 0 0 0 io_in[3]
port 76 nsew signal input
flabel metal3 s 583520 21638 584800 21750 0 FreeSans 1120 0 0 0 io_in[4]
port 77 nsew signal input
flabel metal3 s 583520 48096 584800 48208 0 FreeSans 1120 0 0 0 io_in[5]
port 78 nsew signal input
flabel metal3 s 583520 92754 584800 92866 0 FreeSans 1120 0 0 0 io_in[6]
port 79 nsew signal input
flabel metal3 s 583520 272776 584800 272888 0 FreeSans 1120 0 0 0 io_in[7]
port 80 nsew signal input
flabel metal3 s 583520 317198 584800 317310 0 FreeSans 1120 0 0 0 io_in[8]
port 81 nsew signal input
flabel metal3 s 583520 362420 584800 362532 0 FreeSans 1120 0 0 0 io_in[9]
port 82 nsew signal input
flabel metal3 s 583520 1544 584800 1656 0 FreeSans 1120 0 0 0 io_in_3v3[0]
port 83 nsew signal input
flabel metal3 s 583520 407660 584800 407772 0 FreeSans 1120 0 0 0 io_in_3v3[10]
port 84 nsew signal input
flabel metal3 s 583520 452082 584800 452194 0 FreeSans 1120 0 0 0 io_in_3v3[11]
port 85 nsew signal input
flabel metal3 s 583520 496504 584800 496616 0 FreeSans 1120 0 0 0 io_in_3v3[12]
port 86 nsew signal input
flabel metal3 s 583520 585926 584800 586038 0 FreeSans 1120 0 0 0 io_in_3v3[13]
port 87 nsew signal input
flabel metal3 s -800 509166 480 509278 0 FreeSans 1120 0 0 0 io_in_3v3[14]
port 88 nsew signal input
flabel metal3 s -800 465944 480 466056 0 FreeSans 1120 0 0 0 io_in_3v3[15]
port 89 nsew signal input
flabel metal3 s -800 422722 480 422834 0 FreeSans 1120 0 0 0 io_in_3v3[16]
port 90 nsew signal input
flabel metal3 s -800 379500 480 379612 0 FreeSans 1120 0 0 0 io_in_3v3[17]
port 91 nsew signal input
flabel metal3 s -800 336278 480 336390 0 FreeSans 1120 0 0 0 io_in_3v3[18]
port 92 nsew signal input
flabel metal3 s -800 293056 480 293168 0 FreeSans 1120 0 0 0 io_in_3v3[19]
port 93 nsew signal input
flabel metal3 s 583520 6272 584800 6384 0 FreeSans 1120 0 0 0 io_in_3v3[1]
port 94 nsew signal input
flabel metal3 s -800 250034 480 250146 0 FreeSans 1120 0 0 0 io_in_3v3[20]
port 95 nsew signal input
flabel metal3 s -800 122412 480 122524 0 FreeSans 1120 0 0 0 io_in_3v3[21]
port 96 nsew signal input
flabel metal3 s -800 79190 480 79302 0 FreeSans 1120 0 0 0 io_in_3v3[22]
port 97 nsew signal input
flabel metal3 s -800 35968 480 36080 0 FreeSans 1120 0 0 0 io_in_3v3[23]
port 98 nsew signal input
flabel metal3 s -800 14546 480 14658 0 FreeSans 1120 0 0 0 io_in_3v3[24]
port 99 nsew signal input
flabel metal3 s -800 9818 480 9930 0 FreeSans 1120 0 0 0 io_in_3v3[25]
port 100 nsew signal input
flabel metal3 s -800 5090 480 5202 0 FreeSans 1120 0 0 0 io_in_3v3[26]
port 101 nsew signal input
flabel metal3 s 583520 11000 584800 11112 0 FreeSans 1120 0 0 0 io_in_3v3[2]
port 102 nsew signal input
flabel metal3 s 583520 15728 584800 15840 0 FreeSans 1120 0 0 0 io_in_3v3[3]
port 103 nsew signal input
flabel metal3 s 583520 20456 584800 20568 0 FreeSans 1120 0 0 0 io_in_3v3[4]
port 104 nsew signal input
flabel metal3 s 583520 46914 584800 47026 0 FreeSans 1120 0 0 0 io_in_3v3[5]
port 105 nsew signal input
flabel metal3 s 583520 91572 584800 91684 0 FreeSans 1120 0 0 0 io_in_3v3[6]
port 106 nsew signal input
flabel metal3 s 583520 271594 584800 271706 0 FreeSans 1120 0 0 0 io_in_3v3[7]
port 107 nsew signal input
flabel metal3 s 583520 316016 584800 316128 0 FreeSans 1120 0 0 0 io_in_3v3[8]
port 108 nsew signal input
flabel metal3 s 583520 361238 584800 361350 0 FreeSans 1120 0 0 0 io_in_3v3[9]
port 109 nsew signal input
flabel metal3 s 583520 5090 584800 5202 0 FreeSans 1120 0 0 0 io_oeb[0]
port 110 nsew signal tristate
flabel metal3 s 583520 411206 584800 411318 0 FreeSans 1120 0 0 0 io_oeb[10]
port 111 nsew signal tristate
flabel metal3 s 583520 455628 584800 455740 0 FreeSans 1120 0 0 0 io_oeb[11]
port 112 nsew signal tristate
flabel metal3 s 583520 500050 584800 500162 0 FreeSans 1120 0 0 0 io_oeb[12]
port 113 nsew signal tristate
flabel metal3 s 583520 589472 584800 589584 0 FreeSans 1120 0 0 0 io_oeb[13]
port 114 nsew signal tristate
flabel metal3 s -800 505620 480 505732 0 FreeSans 1120 0 0 0 io_oeb[14]
port 115 nsew signal tristate
flabel metal3 s -800 462398 480 462510 0 FreeSans 1120 0 0 0 io_oeb[15]
port 116 nsew signal tristate
flabel metal3 s -800 419176 480 419288 0 FreeSans 1120 0 0 0 io_oeb[16]
port 117 nsew signal tristate
flabel metal3 s -800 375954 480 376066 0 FreeSans 1120 0 0 0 io_oeb[17]
port 118 nsew signal tristate
flabel metal3 s -800 332732 480 332844 0 FreeSans 1120 0 0 0 io_oeb[18]
port 119 nsew signal tristate
flabel metal3 s -800 289510 480 289622 0 FreeSans 1120 0 0 0 io_oeb[19]
port 120 nsew signal tristate
flabel metal3 s 583520 9818 584800 9930 0 FreeSans 1120 0 0 0 io_oeb[1]
port 121 nsew signal tristate
flabel metal3 s -800 246488 480 246600 0 FreeSans 1120 0 0 0 io_oeb[20]
port 122 nsew signal tristate
flabel metal3 s -800 118866 480 118978 0 FreeSans 1120 0 0 0 io_oeb[21]
port 123 nsew signal tristate
flabel metal3 s -800 75644 480 75756 0 FreeSans 1120 0 0 0 io_oeb[22]
port 124 nsew signal tristate
flabel metal3 s -800 32422 480 32534 0 FreeSans 1120 0 0 0 io_oeb[23]
port 125 nsew signal tristate
flabel metal3 s -800 11000 480 11112 0 FreeSans 1120 0 0 0 io_oeb[24]
port 126 nsew signal tristate
flabel metal3 s -800 6272 480 6384 0 FreeSans 1120 0 0 0 io_oeb[25]
port 127 nsew signal tristate
flabel metal3 s -800 1544 480 1656 0 FreeSans 1120 0 0 0 io_oeb[26]
port 128 nsew signal tristate
flabel metal3 s 583520 14546 584800 14658 0 FreeSans 1120 0 0 0 io_oeb[2]
port 129 nsew signal tristate
flabel metal3 s 583520 19274 584800 19386 0 FreeSans 1120 0 0 0 io_oeb[3]
port 130 nsew signal tristate
flabel metal3 s 583520 24002 584800 24114 0 FreeSans 1120 0 0 0 io_oeb[4]
port 131 nsew signal tristate
flabel metal3 s 583520 50460 584800 50572 0 FreeSans 1120 0 0 0 io_oeb[5]
port 132 nsew signal tristate
flabel metal3 s 583520 95118 584800 95230 0 FreeSans 1120 0 0 0 io_oeb[6]
port 133 nsew signal tristate
flabel metal3 s 583520 275140 584800 275252 0 FreeSans 1120 0 0 0 io_oeb[7]
port 134 nsew signal tristate
flabel metal3 s 583520 319562 584800 319674 0 FreeSans 1120 0 0 0 io_oeb[8]
port 135 nsew signal tristate
flabel metal3 s 583520 364784 584800 364896 0 FreeSans 1120 0 0 0 io_oeb[9]
port 136 nsew signal tristate
flabel metal3 s 583520 3908 584800 4020 0 FreeSans 1120 0 0 0 io_out[0]
port 137 nsew signal tristate
flabel metal3 s 583520 410024 584800 410136 0 FreeSans 1120 0 0 0 io_out[10]
port 138 nsew signal tristate
flabel metal3 s 583520 454446 584800 454558 0 FreeSans 1120 0 0 0 io_out[11]
port 139 nsew signal tristate
flabel metal3 s 583520 498868 584800 498980 0 FreeSans 1120 0 0 0 io_out[12]
port 140 nsew signal tristate
flabel metal3 s 583520 588290 584800 588402 0 FreeSans 1120 0 0 0 io_out[13]
port 141 nsew signal tristate
flabel metal3 s -800 506802 480 506914 0 FreeSans 1120 0 0 0 io_out[14]
port 142 nsew signal tristate
flabel metal3 s -800 463580 480 463692 0 FreeSans 1120 0 0 0 io_out[15]
port 143 nsew signal tristate
flabel metal3 s -800 420358 480 420470 0 FreeSans 1120 0 0 0 io_out[16]
port 144 nsew signal tristate
flabel metal3 s -800 377136 480 377248 0 FreeSans 1120 0 0 0 io_out[17]
port 145 nsew signal tristate
flabel metal3 s -800 333914 480 334026 0 FreeSans 1120 0 0 0 io_out[18]
port 146 nsew signal tristate
flabel metal3 s -800 290692 480 290804 0 FreeSans 1120 0 0 0 io_out[19]
port 147 nsew signal tristate
flabel metal3 s 583520 8636 584800 8748 0 FreeSans 1120 0 0 0 io_out[1]
port 148 nsew signal tristate
flabel metal3 s -800 247670 480 247782 0 FreeSans 1120 0 0 0 io_out[20]
port 149 nsew signal tristate
flabel metal3 s -800 120048 480 120160 0 FreeSans 1120 0 0 0 io_out[21]
port 150 nsew signal tristate
flabel metal3 s -800 76826 480 76938 0 FreeSans 1120 0 0 0 io_out[22]
port 151 nsew signal tristate
flabel metal3 s -800 33604 480 33716 0 FreeSans 1120 0 0 0 io_out[23]
port 152 nsew signal tristate
flabel metal3 s -800 12182 480 12294 0 FreeSans 1120 0 0 0 io_out[24]
port 153 nsew signal tristate
flabel metal3 s -800 7454 480 7566 0 FreeSans 1120 0 0 0 io_out[25]
port 154 nsew signal tristate
flabel metal3 s -800 2726 480 2838 0 FreeSans 1120 0 0 0 io_out[26]
port 155 nsew signal tristate
flabel metal3 s 583520 13364 584800 13476 0 FreeSans 1120 0 0 0 io_out[2]
port 156 nsew signal tristate
flabel metal3 s 583520 18092 584800 18204 0 FreeSans 1120 0 0 0 io_out[3]
port 157 nsew signal tristate
flabel metal3 s 583520 22820 584800 22932 0 FreeSans 1120 0 0 0 io_out[4]
port 158 nsew signal tristate
flabel metal3 s 583520 49278 584800 49390 0 FreeSans 1120 0 0 0 io_out[5]
port 159 nsew signal tristate
flabel metal3 s 583520 93936 584800 94048 0 FreeSans 1120 0 0 0 io_out[6]
port 160 nsew signal tristate
flabel metal3 s 583520 273958 584800 274070 0 FreeSans 1120 0 0 0 io_out[7]
port 161 nsew signal tristate
flabel metal3 s 583520 318380 584800 318492 0 FreeSans 1120 0 0 0 io_out[8]
port 162 nsew signal tristate
flabel metal3 s 583520 363602 584800 363714 0 FreeSans 1120 0 0 0 io_out[9]
port 163 nsew signal tristate
flabel metal2 s 125816 -800 125928 480 0 FreeSans 1120 90 0 0 la_data_in[0]
port 164 nsew signal input
flabel metal2 s 480416 -800 480528 480 0 FreeSans 1120 90 0 0 la_data_in[100]
port 165 nsew signal input
flabel metal2 s 483962 -800 484074 480 0 FreeSans 1120 90 0 0 la_data_in[101]
port 166 nsew signal input
flabel metal2 s 487508 -800 487620 480 0 FreeSans 1120 90 0 0 la_data_in[102]
port 167 nsew signal input
flabel metal2 s 491054 -800 491166 480 0 FreeSans 1120 90 0 0 la_data_in[103]
port 168 nsew signal input
flabel metal2 s 494600 -800 494712 480 0 FreeSans 1120 90 0 0 la_data_in[104]
port 169 nsew signal input
flabel metal2 s 498146 -800 498258 480 0 FreeSans 1120 90 0 0 la_data_in[105]
port 170 nsew signal input
flabel metal2 s 501692 -800 501804 480 0 FreeSans 1120 90 0 0 la_data_in[106]
port 171 nsew signal input
flabel metal2 s 505238 -800 505350 480 0 FreeSans 1120 90 0 0 la_data_in[107]
port 172 nsew signal input
flabel metal2 s 508784 -800 508896 480 0 FreeSans 1120 90 0 0 la_data_in[108]
port 173 nsew signal input
flabel metal2 s 512330 -800 512442 480 0 FreeSans 1120 90 0 0 la_data_in[109]
port 174 nsew signal input
flabel metal2 s 161276 -800 161388 480 0 FreeSans 1120 90 0 0 la_data_in[10]
port 175 nsew signal input
flabel metal2 s 515876 -800 515988 480 0 FreeSans 1120 90 0 0 la_data_in[110]
port 176 nsew signal input
flabel metal2 s 519422 -800 519534 480 0 FreeSans 1120 90 0 0 la_data_in[111]
port 177 nsew signal input
flabel metal2 s 522968 -800 523080 480 0 FreeSans 1120 90 0 0 la_data_in[112]
port 178 nsew signal input
flabel metal2 s 526514 -800 526626 480 0 FreeSans 1120 90 0 0 la_data_in[113]
port 179 nsew signal input
flabel metal2 s 530060 -800 530172 480 0 FreeSans 1120 90 0 0 la_data_in[114]
port 180 nsew signal input
flabel metal2 s 533606 -800 533718 480 0 FreeSans 1120 90 0 0 la_data_in[115]
port 181 nsew signal input
flabel metal2 s 537152 -800 537264 480 0 FreeSans 1120 90 0 0 la_data_in[116]
port 182 nsew signal input
flabel metal2 s 540698 -800 540810 480 0 FreeSans 1120 90 0 0 la_data_in[117]
port 183 nsew signal input
flabel metal2 s 544244 -800 544356 480 0 FreeSans 1120 90 0 0 la_data_in[118]
port 184 nsew signal input
flabel metal2 s 547790 -800 547902 480 0 FreeSans 1120 90 0 0 la_data_in[119]
port 185 nsew signal input
flabel metal2 s 164822 -800 164934 480 0 FreeSans 1120 90 0 0 la_data_in[11]
port 186 nsew signal input
flabel metal2 s 551336 -800 551448 480 0 FreeSans 1120 90 0 0 la_data_in[120]
port 187 nsew signal input
flabel metal2 s 554882 -800 554994 480 0 FreeSans 1120 90 0 0 la_data_in[121]
port 188 nsew signal input
flabel metal2 s 558428 -800 558540 480 0 FreeSans 1120 90 0 0 la_data_in[122]
port 189 nsew signal input
flabel metal2 s 561974 -800 562086 480 0 FreeSans 1120 90 0 0 la_data_in[123]
port 190 nsew signal input
flabel metal2 s 565520 -800 565632 480 0 FreeSans 1120 90 0 0 la_data_in[124]
port 191 nsew signal input
flabel metal2 s 569066 -800 569178 480 0 FreeSans 1120 90 0 0 la_data_in[125]
port 192 nsew signal input
flabel metal2 s 572612 -800 572724 480 0 FreeSans 1120 90 0 0 la_data_in[126]
port 193 nsew signal input
flabel metal2 s 576158 -800 576270 480 0 FreeSans 1120 90 0 0 la_data_in[127]
port 194 nsew signal input
flabel metal2 s 168368 -800 168480 480 0 FreeSans 1120 90 0 0 la_data_in[12]
port 195 nsew signal input
flabel metal2 s 171914 -800 172026 480 0 FreeSans 1120 90 0 0 la_data_in[13]
port 196 nsew signal input
flabel metal2 s 175460 -800 175572 480 0 FreeSans 1120 90 0 0 la_data_in[14]
port 197 nsew signal input
flabel metal2 s 179006 -800 179118 480 0 FreeSans 1120 90 0 0 la_data_in[15]
port 198 nsew signal input
flabel metal2 s 182552 -800 182664 480 0 FreeSans 1120 90 0 0 la_data_in[16]
port 199 nsew signal input
flabel metal2 s 186098 -800 186210 480 0 FreeSans 1120 90 0 0 la_data_in[17]
port 200 nsew signal input
flabel metal2 s 189644 -800 189756 480 0 FreeSans 1120 90 0 0 la_data_in[18]
port 201 nsew signal input
flabel metal2 s 193190 -800 193302 480 0 FreeSans 1120 90 0 0 la_data_in[19]
port 202 nsew signal input
flabel metal2 s 129362 -800 129474 480 0 FreeSans 1120 90 0 0 la_data_in[1]
port 203 nsew signal input
flabel metal2 s 196736 -800 196848 480 0 FreeSans 1120 90 0 0 la_data_in[20]
port 204 nsew signal input
flabel metal2 s 200282 -800 200394 480 0 FreeSans 1120 90 0 0 la_data_in[21]
port 205 nsew signal input
flabel metal2 s 203828 -800 203940 480 0 FreeSans 1120 90 0 0 la_data_in[22]
port 206 nsew signal input
flabel metal2 s 207374 -800 207486 480 0 FreeSans 1120 90 0 0 la_data_in[23]
port 207 nsew signal input
flabel metal2 s 210920 -800 211032 480 0 FreeSans 1120 90 0 0 la_data_in[24]
port 208 nsew signal input
flabel metal2 s 214466 -800 214578 480 0 FreeSans 1120 90 0 0 la_data_in[25]
port 209 nsew signal input
flabel metal2 s 218012 -800 218124 480 0 FreeSans 1120 90 0 0 la_data_in[26]
port 210 nsew signal input
flabel metal2 s 221558 -800 221670 480 0 FreeSans 1120 90 0 0 la_data_in[27]
port 211 nsew signal input
flabel metal2 s 225104 -800 225216 480 0 FreeSans 1120 90 0 0 la_data_in[28]
port 212 nsew signal input
flabel metal2 s 228650 -800 228762 480 0 FreeSans 1120 90 0 0 la_data_in[29]
port 213 nsew signal input
flabel metal2 s 132908 -800 133020 480 0 FreeSans 1120 90 0 0 la_data_in[2]
port 214 nsew signal input
flabel metal2 s 232196 -800 232308 480 0 FreeSans 1120 90 0 0 la_data_in[30]
port 215 nsew signal input
flabel metal2 s 235742 -800 235854 480 0 FreeSans 1120 90 0 0 la_data_in[31]
port 216 nsew signal input
flabel metal2 s 239288 -800 239400 480 0 FreeSans 1120 90 0 0 la_data_in[32]
port 217 nsew signal input
flabel metal2 s 242834 -800 242946 480 0 FreeSans 1120 90 0 0 la_data_in[33]
port 218 nsew signal input
flabel metal2 s 246380 -800 246492 480 0 FreeSans 1120 90 0 0 la_data_in[34]
port 219 nsew signal input
flabel metal2 s 249926 -800 250038 480 0 FreeSans 1120 90 0 0 la_data_in[35]
port 220 nsew signal input
flabel metal2 s 253472 -800 253584 480 0 FreeSans 1120 90 0 0 la_data_in[36]
port 221 nsew signal input
flabel metal2 s 257018 -800 257130 480 0 FreeSans 1120 90 0 0 la_data_in[37]
port 222 nsew signal input
flabel metal2 s 260564 -800 260676 480 0 FreeSans 1120 90 0 0 la_data_in[38]
port 223 nsew signal input
flabel metal2 s 264110 -800 264222 480 0 FreeSans 1120 90 0 0 la_data_in[39]
port 224 nsew signal input
flabel metal2 s 136454 -800 136566 480 0 FreeSans 1120 90 0 0 la_data_in[3]
port 225 nsew signal input
flabel metal2 s 267656 -800 267768 480 0 FreeSans 1120 90 0 0 la_data_in[40]
port 226 nsew signal input
flabel metal2 s 271202 -800 271314 480 0 FreeSans 1120 90 0 0 la_data_in[41]
port 227 nsew signal input
flabel metal2 s 274748 -800 274860 480 0 FreeSans 1120 90 0 0 la_data_in[42]
port 228 nsew signal input
flabel metal2 s 278294 -800 278406 480 0 FreeSans 1120 90 0 0 la_data_in[43]
port 229 nsew signal input
flabel metal2 s 281840 -800 281952 480 0 FreeSans 1120 90 0 0 la_data_in[44]
port 230 nsew signal input
flabel metal2 s 285386 -800 285498 480 0 FreeSans 1120 90 0 0 la_data_in[45]
port 231 nsew signal input
flabel metal2 s 288932 -800 289044 480 0 FreeSans 1120 90 0 0 la_data_in[46]
port 232 nsew signal input
flabel metal2 s 292478 -800 292590 480 0 FreeSans 1120 90 0 0 la_data_in[47]
port 233 nsew signal input
flabel metal2 s 296024 -800 296136 480 0 FreeSans 1120 90 0 0 la_data_in[48]
port 234 nsew signal input
flabel metal2 s 299570 -800 299682 480 0 FreeSans 1120 90 0 0 la_data_in[49]
port 235 nsew signal input
flabel metal2 s 140000 -800 140112 480 0 FreeSans 1120 90 0 0 la_data_in[4]
port 236 nsew signal input
flabel metal2 s 303116 -800 303228 480 0 FreeSans 1120 90 0 0 la_data_in[50]
port 237 nsew signal input
flabel metal2 s 306662 -800 306774 480 0 FreeSans 1120 90 0 0 la_data_in[51]
port 238 nsew signal input
flabel metal2 s 310208 -800 310320 480 0 FreeSans 1120 90 0 0 la_data_in[52]
port 239 nsew signal input
flabel metal2 s 313754 -800 313866 480 0 FreeSans 1120 90 0 0 la_data_in[53]
port 240 nsew signal input
flabel metal2 s 317300 -800 317412 480 0 FreeSans 1120 90 0 0 la_data_in[54]
port 241 nsew signal input
flabel metal2 s 320846 -800 320958 480 0 FreeSans 1120 90 0 0 la_data_in[55]
port 242 nsew signal input
flabel metal2 s 324392 -800 324504 480 0 FreeSans 1120 90 0 0 la_data_in[56]
port 243 nsew signal input
flabel metal2 s 327938 -800 328050 480 0 FreeSans 1120 90 0 0 la_data_in[57]
port 244 nsew signal input
flabel metal2 s 331484 -800 331596 480 0 FreeSans 1120 90 0 0 la_data_in[58]
port 245 nsew signal input
flabel metal2 s 335030 -800 335142 480 0 FreeSans 1120 90 0 0 la_data_in[59]
port 246 nsew signal input
flabel metal2 s 143546 -800 143658 480 0 FreeSans 1120 90 0 0 la_data_in[5]
port 247 nsew signal input
flabel metal2 s 338576 -800 338688 480 0 FreeSans 1120 90 0 0 la_data_in[60]
port 248 nsew signal input
flabel metal2 s 342122 -800 342234 480 0 FreeSans 1120 90 0 0 la_data_in[61]
port 249 nsew signal input
flabel metal2 s 345668 -800 345780 480 0 FreeSans 1120 90 0 0 la_data_in[62]
port 250 nsew signal input
flabel metal2 s 349214 -800 349326 480 0 FreeSans 1120 90 0 0 la_data_in[63]
port 251 nsew signal input
flabel metal2 s 352760 -800 352872 480 0 FreeSans 1120 90 0 0 la_data_in[64]
port 252 nsew signal input
flabel metal2 s 356306 -800 356418 480 0 FreeSans 1120 90 0 0 la_data_in[65]
port 253 nsew signal input
flabel metal2 s 359852 -800 359964 480 0 FreeSans 1120 90 0 0 la_data_in[66]
port 254 nsew signal input
flabel metal2 s 363398 -800 363510 480 0 FreeSans 1120 90 0 0 la_data_in[67]
port 255 nsew signal input
flabel metal2 s 366944 -800 367056 480 0 FreeSans 1120 90 0 0 la_data_in[68]
port 256 nsew signal input
flabel metal2 s 370490 -800 370602 480 0 FreeSans 1120 90 0 0 la_data_in[69]
port 257 nsew signal input
flabel metal2 s 147092 -800 147204 480 0 FreeSans 1120 90 0 0 la_data_in[6]
port 258 nsew signal input
flabel metal2 s 374036 -800 374148 480 0 FreeSans 1120 90 0 0 la_data_in[70]
port 259 nsew signal input
flabel metal2 s 377582 -800 377694 480 0 FreeSans 1120 90 0 0 la_data_in[71]
port 260 nsew signal input
flabel metal2 s 381128 -800 381240 480 0 FreeSans 1120 90 0 0 la_data_in[72]
port 261 nsew signal input
flabel metal2 s 384674 -800 384786 480 0 FreeSans 1120 90 0 0 la_data_in[73]
port 262 nsew signal input
flabel metal2 s 388220 -800 388332 480 0 FreeSans 1120 90 0 0 la_data_in[74]
port 263 nsew signal input
flabel metal2 s 391766 -800 391878 480 0 FreeSans 1120 90 0 0 la_data_in[75]
port 264 nsew signal input
flabel metal2 s 395312 -800 395424 480 0 FreeSans 1120 90 0 0 la_data_in[76]
port 265 nsew signal input
flabel metal2 s 398858 -800 398970 480 0 FreeSans 1120 90 0 0 la_data_in[77]
port 266 nsew signal input
flabel metal2 s 402404 -800 402516 480 0 FreeSans 1120 90 0 0 la_data_in[78]
port 267 nsew signal input
flabel metal2 s 405950 -800 406062 480 0 FreeSans 1120 90 0 0 la_data_in[79]
port 268 nsew signal input
flabel metal2 s 150638 -800 150750 480 0 FreeSans 1120 90 0 0 la_data_in[7]
port 269 nsew signal input
flabel metal2 s 409496 -800 409608 480 0 FreeSans 1120 90 0 0 la_data_in[80]
port 270 nsew signal input
flabel metal2 s 413042 -800 413154 480 0 FreeSans 1120 90 0 0 la_data_in[81]
port 271 nsew signal input
flabel metal2 s 416588 -800 416700 480 0 FreeSans 1120 90 0 0 la_data_in[82]
port 272 nsew signal input
flabel metal2 s 420134 -800 420246 480 0 FreeSans 1120 90 0 0 la_data_in[83]
port 273 nsew signal input
flabel metal2 s 423680 -800 423792 480 0 FreeSans 1120 90 0 0 la_data_in[84]
port 274 nsew signal input
flabel metal2 s 427226 -800 427338 480 0 FreeSans 1120 90 0 0 la_data_in[85]
port 275 nsew signal input
flabel metal2 s 430772 -800 430884 480 0 FreeSans 1120 90 0 0 la_data_in[86]
port 276 nsew signal input
flabel metal2 s 434318 -800 434430 480 0 FreeSans 1120 90 0 0 la_data_in[87]
port 277 nsew signal input
flabel metal2 s 437864 -800 437976 480 0 FreeSans 1120 90 0 0 la_data_in[88]
port 278 nsew signal input
flabel metal2 s 441410 -800 441522 480 0 FreeSans 1120 90 0 0 la_data_in[89]
port 279 nsew signal input
flabel metal2 s 154184 -800 154296 480 0 FreeSans 1120 90 0 0 la_data_in[8]
port 280 nsew signal input
flabel metal2 s 444956 -800 445068 480 0 FreeSans 1120 90 0 0 la_data_in[90]
port 281 nsew signal input
flabel metal2 s 448502 -800 448614 480 0 FreeSans 1120 90 0 0 la_data_in[91]
port 282 nsew signal input
flabel metal2 s 452048 -800 452160 480 0 FreeSans 1120 90 0 0 la_data_in[92]
port 283 nsew signal input
flabel metal2 s 455594 -800 455706 480 0 FreeSans 1120 90 0 0 la_data_in[93]
port 284 nsew signal input
flabel metal2 s 459140 -800 459252 480 0 FreeSans 1120 90 0 0 la_data_in[94]
port 285 nsew signal input
flabel metal2 s 462686 -800 462798 480 0 FreeSans 1120 90 0 0 la_data_in[95]
port 286 nsew signal input
flabel metal2 s 466232 -800 466344 480 0 FreeSans 1120 90 0 0 la_data_in[96]
port 287 nsew signal input
flabel metal2 s 469778 -800 469890 480 0 FreeSans 1120 90 0 0 la_data_in[97]
port 288 nsew signal input
flabel metal2 s 473324 -800 473436 480 0 FreeSans 1120 90 0 0 la_data_in[98]
port 289 nsew signal input
flabel metal2 s 476870 -800 476982 480 0 FreeSans 1120 90 0 0 la_data_in[99]
port 290 nsew signal input
flabel metal2 s 157730 -800 157842 480 0 FreeSans 1120 90 0 0 la_data_in[9]
port 291 nsew signal input
flabel metal2 s 126998 -800 127110 480 0 FreeSans 1120 90 0 0 la_data_out[0]
port 292 nsew signal tristate
flabel metal2 s 481598 -800 481710 480 0 FreeSans 1120 90 0 0 la_data_out[100]
port 293 nsew signal tristate
flabel metal2 s 485144 -800 485256 480 0 FreeSans 1120 90 0 0 la_data_out[101]
port 294 nsew signal tristate
flabel metal2 s 488690 -800 488802 480 0 FreeSans 1120 90 0 0 la_data_out[102]
port 295 nsew signal tristate
flabel metal2 s 492236 -800 492348 480 0 FreeSans 1120 90 0 0 la_data_out[103]
port 296 nsew signal tristate
flabel metal2 s 495782 -800 495894 480 0 FreeSans 1120 90 0 0 la_data_out[104]
port 297 nsew signal tristate
flabel metal2 s 499328 -800 499440 480 0 FreeSans 1120 90 0 0 la_data_out[105]
port 298 nsew signal tristate
flabel metal2 s 502874 -800 502986 480 0 FreeSans 1120 90 0 0 la_data_out[106]
port 299 nsew signal tristate
flabel metal2 s 506420 -800 506532 480 0 FreeSans 1120 90 0 0 la_data_out[107]
port 300 nsew signal tristate
flabel metal2 s 509966 -800 510078 480 0 FreeSans 1120 90 0 0 la_data_out[108]
port 301 nsew signal tristate
flabel metal2 s 513512 -800 513624 480 0 FreeSans 1120 90 0 0 la_data_out[109]
port 302 nsew signal tristate
flabel metal2 s 162458 -800 162570 480 0 FreeSans 1120 90 0 0 la_data_out[10]
port 303 nsew signal tristate
flabel metal2 s 517058 -800 517170 480 0 FreeSans 1120 90 0 0 la_data_out[110]
port 304 nsew signal tristate
flabel metal2 s 520604 -800 520716 480 0 FreeSans 1120 90 0 0 la_data_out[111]
port 305 nsew signal tristate
flabel metal2 s 524150 -800 524262 480 0 FreeSans 1120 90 0 0 la_data_out[112]
port 306 nsew signal tristate
flabel metal2 s 527696 -800 527808 480 0 FreeSans 1120 90 0 0 la_data_out[113]
port 307 nsew signal tristate
flabel metal2 s 531242 -800 531354 480 0 FreeSans 1120 90 0 0 la_data_out[114]
port 308 nsew signal tristate
flabel metal2 s 534788 -800 534900 480 0 FreeSans 1120 90 0 0 la_data_out[115]
port 309 nsew signal tristate
flabel metal2 s 538334 -800 538446 480 0 FreeSans 1120 90 0 0 la_data_out[116]
port 310 nsew signal tristate
flabel metal2 s 541880 -800 541992 480 0 FreeSans 1120 90 0 0 la_data_out[117]
port 311 nsew signal tristate
flabel metal2 s 545426 -800 545538 480 0 FreeSans 1120 90 0 0 la_data_out[118]
port 312 nsew signal tristate
flabel metal2 s 548972 -800 549084 480 0 FreeSans 1120 90 0 0 la_data_out[119]
port 313 nsew signal tristate
flabel metal2 s 166004 -800 166116 480 0 FreeSans 1120 90 0 0 la_data_out[11]
port 314 nsew signal tristate
flabel metal2 s 552518 -800 552630 480 0 FreeSans 1120 90 0 0 la_data_out[120]
port 315 nsew signal tristate
flabel metal2 s 556064 -800 556176 480 0 FreeSans 1120 90 0 0 la_data_out[121]
port 316 nsew signal tristate
flabel metal2 s 559610 -800 559722 480 0 FreeSans 1120 90 0 0 la_data_out[122]
port 317 nsew signal tristate
flabel metal2 s 563156 -800 563268 480 0 FreeSans 1120 90 0 0 la_data_out[123]
port 318 nsew signal tristate
flabel metal2 s 566702 -800 566814 480 0 FreeSans 1120 90 0 0 la_data_out[124]
port 319 nsew signal tristate
flabel metal2 s 570248 -800 570360 480 0 FreeSans 1120 90 0 0 la_data_out[125]
port 320 nsew signal tristate
flabel metal2 s 573794 -800 573906 480 0 FreeSans 1120 90 0 0 la_data_out[126]
port 321 nsew signal tristate
flabel metal2 s 577340 -800 577452 480 0 FreeSans 1120 90 0 0 la_data_out[127]
port 322 nsew signal tristate
flabel metal2 s 169550 -800 169662 480 0 FreeSans 1120 90 0 0 la_data_out[12]
port 323 nsew signal tristate
flabel metal2 s 173096 -800 173208 480 0 FreeSans 1120 90 0 0 la_data_out[13]
port 324 nsew signal tristate
flabel metal2 s 176642 -800 176754 480 0 FreeSans 1120 90 0 0 la_data_out[14]
port 325 nsew signal tristate
flabel metal2 s 180188 -800 180300 480 0 FreeSans 1120 90 0 0 la_data_out[15]
port 326 nsew signal tristate
flabel metal2 s 183734 -800 183846 480 0 FreeSans 1120 90 0 0 la_data_out[16]
port 327 nsew signal tristate
flabel metal2 s 187280 -800 187392 480 0 FreeSans 1120 90 0 0 la_data_out[17]
port 328 nsew signal tristate
flabel metal2 s 190826 -800 190938 480 0 FreeSans 1120 90 0 0 la_data_out[18]
port 329 nsew signal tristate
flabel metal2 s 194372 -800 194484 480 0 FreeSans 1120 90 0 0 la_data_out[19]
port 330 nsew signal tristate
flabel metal2 s 130544 -800 130656 480 0 FreeSans 1120 90 0 0 la_data_out[1]
port 331 nsew signal tristate
flabel metal2 s 197918 -800 198030 480 0 FreeSans 1120 90 0 0 la_data_out[20]
port 332 nsew signal tristate
flabel metal2 s 201464 -800 201576 480 0 FreeSans 1120 90 0 0 la_data_out[21]
port 333 nsew signal tristate
flabel metal2 s 205010 -800 205122 480 0 FreeSans 1120 90 0 0 la_data_out[22]
port 334 nsew signal tristate
flabel metal2 s 208556 -800 208668 480 0 FreeSans 1120 90 0 0 la_data_out[23]
port 335 nsew signal tristate
flabel metal2 s 212102 -800 212214 480 0 FreeSans 1120 90 0 0 la_data_out[24]
port 336 nsew signal tristate
flabel metal2 s 215648 -800 215760 480 0 FreeSans 1120 90 0 0 la_data_out[25]
port 337 nsew signal tristate
flabel metal2 s 219194 -800 219306 480 0 FreeSans 1120 90 0 0 la_data_out[26]
port 338 nsew signal tristate
flabel metal2 s 222740 -800 222852 480 0 FreeSans 1120 90 0 0 la_data_out[27]
port 339 nsew signal tristate
flabel metal2 s 226286 -800 226398 480 0 FreeSans 1120 90 0 0 la_data_out[28]
port 340 nsew signal tristate
flabel metal2 s 229832 -800 229944 480 0 FreeSans 1120 90 0 0 la_data_out[29]
port 341 nsew signal tristate
flabel metal2 s 134090 -800 134202 480 0 FreeSans 1120 90 0 0 la_data_out[2]
port 342 nsew signal tristate
flabel metal2 s 233378 -800 233490 480 0 FreeSans 1120 90 0 0 la_data_out[30]
port 343 nsew signal tristate
flabel metal2 s 236924 -800 237036 480 0 FreeSans 1120 90 0 0 la_data_out[31]
port 344 nsew signal tristate
flabel metal2 s 240470 -800 240582 480 0 FreeSans 1120 90 0 0 la_data_out[32]
port 345 nsew signal tristate
flabel metal2 s 244016 -800 244128 480 0 FreeSans 1120 90 0 0 la_data_out[33]
port 346 nsew signal tristate
flabel metal2 s 247562 -800 247674 480 0 FreeSans 1120 90 0 0 la_data_out[34]
port 347 nsew signal tristate
flabel metal2 s 251108 -800 251220 480 0 FreeSans 1120 90 0 0 la_data_out[35]
port 348 nsew signal tristate
flabel metal2 s 254654 -800 254766 480 0 FreeSans 1120 90 0 0 la_data_out[36]
port 349 nsew signal tristate
flabel metal2 s 258200 -800 258312 480 0 FreeSans 1120 90 0 0 la_data_out[37]
port 350 nsew signal tristate
flabel metal2 s 261746 -800 261858 480 0 FreeSans 1120 90 0 0 la_data_out[38]
port 351 nsew signal tristate
flabel metal2 s 265292 -800 265404 480 0 FreeSans 1120 90 0 0 la_data_out[39]
port 352 nsew signal tristate
flabel metal2 s 137636 -800 137748 480 0 FreeSans 1120 90 0 0 la_data_out[3]
port 353 nsew signal tristate
flabel metal2 s 268838 -800 268950 480 0 FreeSans 1120 90 0 0 la_data_out[40]
port 354 nsew signal tristate
flabel metal2 s 272384 -800 272496 480 0 FreeSans 1120 90 0 0 la_data_out[41]
port 355 nsew signal tristate
flabel metal2 s 275930 -800 276042 480 0 FreeSans 1120 90 0 0 la_data_out[42]
port 356 nsew signal tristate
flabel metal2 s 279476 -800 279588 480 0 FreeSans 1120 90 0 0 la_data_out[43]
port 357 nsew signal tristate
flabel metal2 s 283022 -800 283134 480 0 FreeSans 1120 90 0 0 la_data_out[44]
port 358 nsew signal tristate
flabel metal2 s 286568 -800 286680 480 0 FreeSans 1120 90 0 0 la_data_out[45]
port 359 nsew signal tristate
flabel metal2 s 290114 -800 290226 480 0 FreeSans 1120 90 0 0 la_data_out[46]
port 360 nsew signal tristate
flabel metal2 s 293660 -800 293772 480 0 FreeSans 1120 90 0 0 la_data_out[47]
port 361 nsew signal tristate
flabel metal2 s 297206 -800 297318 480 0 FreeSans 1120 90 0 0 la_data_out[48]
port 362 nsew signal tristate
flabel metal2 s 300752 -800 300864 480 0 FreeSans 1120 90 0 0 la_data_out[49]
port 363 nsew signal tristate
flabel metal2 s 141182 -800 141294 480 0 FreeSans 1120 90 0 0 la_data_out[4]
port 364 nsew signal tristate
flabel metal2 s 304298 -800 304410 480 0 FreeSans 1120 90 0 0 la_data_out[50]
port 365 nsew signal tristate
flabel metal2 s 307844 -800 307956 480 0 FreeSans 1120 90 0 0 la_data_out[51]
port 366 nsew signal tristate
flabel metal2 s 311390 -800 311502 480 0 FreeSans 1120 90 0 0 la_data_out[52]
port 367 nsew signal tristate
flabel metal2 s 314936 -800 315048 480 0 FreeSans 1120 90 0 0 la_data_out[53]
port 368 nsew signal tristate
flabel metal2 s 318482 -800 318594 480 0 FreeSans 1120 90 0 0 la_data_out[54]
port 369 nsew signal tristate
flabel metal2 s 322028 -800 322140 480 0 FreeSans 1120 90 0 0 la_data_out[55]
port 370 nsew signal tristate
flabel metal2 s 325574 -800 325686 480 0 FreeSans 1120 90 0 0 la_data_out[56]
port 371 nsew signal tristate
flabel metal2 s 329120 -800 329232 480 0 FreeSans 1120 90 0 0 la_data_out[57]
port 372 nsew signal tristate
flabel metal2 s 332666 -800 332778 480 0 FreeSans 1120 90 0 0 la_data_out[58]
port 373 nsew signal tristate
flabel metal2 s 336212 -800 336324 480 0 FreeSans 1120 90 0 0 la_data_out[59]
port 374 nsew signal tristate
flabel metal2 s 144728 -800 144840 480 0 FreeSans 1120 90 0 0 la_data_out[5]
port 375 nsew signal tristate
flabel metal2 s 339758 -800 339870 480 0 FreeSans 1120 90 0 0 la_data_out[60]
port 376 nsew signal tristate
flabel metal2 s 343304 -800 343416 480 0 FreeSans 1120 90 0 0 la_data_out[61]
port 377 nsew signal tristate
flabel metal2 s 346850 -800 346962 480 0 FreeSans 1120 90 0 0 la_data_out[62]
port 378 nsew signal tristate
flabel metal2 s 350396 -800 350508 480 0 FreeSans 1120 90 0 0 la_data_out[63]
port 379 nsew signal tristate
flabel metal2 s 353942 -800 354054 480 0 FreeSans 1120 90 0 0 la_data_out[64]
port 380 nsew signal tristate
flabel metal2 s 357488 -800 357600 480 0 FreeSans 1120 90 0 0 la_data_out[65]
port 381 nsew signal tristate
flabel metal2 s 361034 -800 361146 480 0 FreeSans 1120 90 0 0 la_data_out[66]
port 382 nsew signal tristate
flabel metal2 s 364580 -800 364692 480 0 FreeSans 1120 90 0 0 la_data_out[67]
port 383 nsew signal tristate
flabel metal2 s 368126 -800 368238 480 0 FreeSans 1120 90 0 0 la_data_out[68]
port 384 nsew signal tristate
flabel metal2 s 371672 -800 371784 480 0 FreeSans 1120 90 0 0 la_data_out[69]
port 385 nsew signal tristate
flabel metal2 s 148274 -800 148386 480 0 FreeSans 1120 90 0 0 la_data_out[6]
port 386 nsew signal tristate
flabel metal2 s 375218 -800 375330 480 0 FreeSans 1120 90 0 0 la_data_out[70]
port 387 nsew signal tristate
flabel metal2 s 378764 -800 378876 480 0 FreeSans 1120 90 0 0 la_data_out[71]
port 388 nsew signal tristate
flabel metal2 s 382310 -800 382422 480 0 FreeSans 1120 90 0 0 la_data_out[72]
port 389 nsew signal tristate
flabel metal2 s 385856 -800 385968 480 0 FreeSans 1120 90 0 0 la_data_out[73]
port 390 nsew signal tristate
flabel metal2 s 389402 -800 389514 480 0 FreeSans 1120 90 0 0 la_data_out[74]
port 391 nsew signal tristate
flabel metal2 s 392948 -800 393060 480 0 FreeSans 1120 90 0 0 la_data_out[75]
port 392 nsew signal tristate
flabel metal2 s 396494 -800 396606 480 0 FreeSans 1120 90 0 0 la_data_out[76]
port 393 nsew signal tristate
flabel metal2 s 400040 -800 400152 480 0 FreeSans 1120 90 0 0 la_data_out[77]
port 394 nsew signal tristate
flabel metal2 s 403586 -800 403698 480 0 FreeSans 1120 90 0 0 la_data_out[78]
port 395 nsew signal tristate
flabel metal2 s 407132 -800 407244 480 0 FreeSans 1120 90 0 0 la_data_out[79]
port 396 nsew signal tristate
flabel metal2 s 151820 -800 151932 480 0 FreeSans 1120 90 0 0 la_data_out[7]
port 397 nsew signal tristate
flabel metal2 s 410678 -800 410790 480 0 FreeSans 1120 90 0 0 la_data_out[80]
port 398 nsew signal tristate
flabel metal2 s 414224 -800 414336 480 0 FreeSans 1120 90 0 0 la_data_out[81]
port 399 nsew signal tristate
flabel metal2 s 417770 -800 417882 480 0 FreeSans 1120 90 0 0 la_data_out[82]
port 400 nsew signal tristate
flabel metal2 s 421316 -800 421428 480 0 FreeSans 1120 90 0 0 la_data_out[83]
port 401 nsew signal tristate
flabel metal2 s 424862 -800 424974 480 0 FreeSans 1120 90 0 0 la_data_out[84]
port 402 nsew signal tristate
flabel metal2 s 428408 -800 428520 480 0 FreeSans 1120 90 0 0 la_data_out[85]
port 403 nsew signal tristate
flabel metal2 s 431954 -800 432066 480 0 FreeSans 1120 90 0 0 la_data_out[86]
port 404 nsew signal tristate
flabel metal2 s 435500 -800 435612 480 0 FreeSans 1120 90 0 0 la_data_out[87]
port 405 nsew signal tristate
flabel metal2 s 439046 -800 439158 480 0 FreeSans 1120 90 0 0 la_data_out[88]
port 406 nsew signal tristate
flabel metal2 s 442592 -800 442704 480 0 FreeSans 1120 90 0 0 la_data_out[89]
port 407 nsew signal tristate
flabel metal2 s 155366 -800 155478 480 0 FreeSans 1120 90 0 0 la_data_out[8]
port 408 nsew signal tristate
flabel metal2 s 446138 -800 446250 480 0 FreeSans 1120 90 0 0 la_data_out[90]
port 409 nsew signal tristate
flabel metal2 s 449684 -800 449796 480 0 FreeSans 1120 90 0 0 la_data_out[91]
port 410 nsew signal tristate
flabel metal2 s 453230 -800 453342 480 0 FreeSans 1120 90 0 0 la_data_out[92]
port 411 nsew signal tristate
flabel metal2 s 456776 -800 456888 480 0 FreeSans 1120 90 0 0 la_data_out[93]
port 412 nsew signal tristate
flabel metal2 s 460322 -800 460434 480 0 FreeSans 1120 90 0 0 la_data_out[94]
port 413 nsew signal tristate
flabel metal2 s 463868 -800 463980 480 0 FreeSans 1120 90 0 0 la_data_out[95]
port 414 nsew signal tristate
flabel metal2 s 467414 -800 467526 480 0 FreeSans 1120 90 0 0 la_data_out[96]
port 415 nsew signal tristate
flabel metal2 s 470960 -800 471072 480 0 FreeSans 1120 90 0 0 la_data_out[97]
port 416 nsew signal tristate
flabel metal2 s 474506 -800 474618 480 0 FreeSans 1120 90 0 0 la_data_out[98]
port 417 nsew signal tristate
flabel metal2 s 478052 -800 478164 480 0 FreeSans 1120 90 0 0 la_data_out[99]
port 418 nsew signal tristate
flabel metal2 s 158912 -800 159024 480 0 FreeSans 1120 90 0 0 la_data_out[9]
port 419 nsew signal tristate
flabel metal2 s 128180 -800 128292 480 0 FreeSans 1120 90 0 0 la_oenb[0]
port 420 nsew signal input
flabel metal2 s 482780 -800 482892 480 0 FreeSans 1120 90 0 0 la_oenb[100]
port 421 nsew signal input
flabel metal2 s 486326 -800 486438 480 0 FreeSans 1120 90 0 0 la_oenb[101]
port 422 nsew signal input
flabel metal2 s 489872 -800 489984 480 0 FreeSans 1120 90 0 0 la_oenb[102]
port 423 nsew signal input
flabel metal2 s 493418 -800 493530 480 0 FreeSans 1120 90 0 0 la_oenb[103]
port 424 nsew signal input
flabel metal2 s 496964 -800 497076 480 0 FreeSans 1120 90 0 0 la_oenb[104]
port 425 nsew signal input
flabel metal2 s 500510 -800 500622 480 0 FreeSans 1120 90 0 0 la_oenb[105]
port 426 nsew signal input
flabel metal2 s 504056 -800 504168 480 0 FreeSans 1120 90 0 0 la_oenb[106]
port 427 nsew signal input
flabel metal2 s 507602 -800 507714 480 0 FreeSans 1120 90 0 0 la_oenb[107]
port 428 nsew signal input
flabel metal2 s 511148 -800 511260 480 0 FreeSans 1120 90 0 0 la_oenb[108]
port 429 nsew signal input
flabel metal2 s 514694 -800 514806 480 0 FreeSans 1120 90 0 0 la_oenb[109]
port 430 nsew signal input
flabel metal2 s 163640 -800 163752 480 0 FreeSans 1120 90 0 0 la_oenb[10]
port 431 nsew signal input
flabel metal2 s 518240 -800 518352 480 0 FreeSans 1120 90 0 0 la_oenb[110]
port 432 nsew signal input
flabel metal2 s 521786 -800 521898 480 0 FreeSans 1120 90 0 0 la_oenb[111]
port 433 nsew signal input
flabel metal2 s 525332 -800 525444 480 0 FreeSans 1120 90 0 0 la_oenb[112]
port 434 nsew signal input
flabel metal2 s 528878 -800 528990 480 0 FreeSans 1120 90 0 0 la_oenb[113]
port 435 nsew signal input
flabel metal2 s 532424 -800 532536 480 0 FreeSans 1120 90 0 0 la_oenb[114]
port 436 nsew signal input
flabel metal2 s 535970 -800 536082 480 0 FreeSans 1120 90 0 0 la_oenb[115]
port 437 nsew signal input
flabel metal2 s 539516 -800 539628 480 0 FreeSans 1120 90 0 0 la_oenb[116]
port 438 nsew signal input
flabel metal2 s 543062 -800 543174 480 0 FreeSans 1120 90 0 0 la_oenb[117]
port 439 nsew signal input
flabel metal2 s 546608 -800 546720 480 0 FreeSans 1120 90 0 0 la_oenb[118]
port 440 nsew signal input
flabel metal2 s 550154 -800 550266 480 0 FreeSans 1120 90 0 0 la_oenb[119]
port 441 nsew signal input
flabel metal2 s 167186 -800 167298 480 0 FreeSans 1120 90 0 0 la_oenb[11]
port 442 nsew signal input
flabel metal2 s 553700 -800 553812 480 0 FreeSans 1120 90 0 0 la_oenb[120]
port 443 nsew signal input
flabel metal2 s 557246 -800 557358 480 0 FreeSans 1120 90 0 0 la_oenb[121]
port 444 nsew signal input
flabel metal2 s 560792 -800 560904 480 0 FreeSans 1120 90 0 0 la_oenb[122]
port 445 nsew signal input
flabel metal2 s 564338 -800 564450 480 0 FreeSans 1120 90 0 0 la_oenb[123]
port 446 nsew signal input
flabel metal2 s 567884 -800 567996 480 0 FreeSans 1120 90 0 0 la_oenb[124]
port 447 nsew signal input
flabel metal2 s 571430 -800 571542 480 0 FreeSans 1120 90 0 0 la_oenb[125]
port 448 nsew signal input
flabel metal2 s 574976 -800 575088 480 0 FreeSans 1120 90 0 0 la_oenb[126]
port 449 nsew signal input
flabel metal2 s 578522 -800 578634 480 0 FreeSans 1120 90 0 0 la_oenb[127]
port 450 nsew signal input
flabel metal2 s 170732 -800 170844 480 0 FreeSans 1120 90 0 0 la_oenb[12]
port 451 nsew signal input
flabel metal2 s 174278 -800 174390 480 0 FreeSans 1120 90 0 0 la_oenb[13]
port 452 nsew signal input
flabel metal2 s 177824 -800 177936 480 0 FreeSans 1120 90 0 0 la_oenb[14]
port 453 nsew signal input
flabel metal2 s 181370 -800 181482 480 0 FreeSans 1120 90 0 0 la_oenb[15]
port 454 nsew signal input
flabel metal2 s 184916 -800 185028 480 0 FreeSans 1120 90 0 0 la_oenb[16]
port 455 nsew signal input
flabel metal2 s 188462 -800 188574 480 0 FreeSans 1120 90 0 0 la_oenb[17]
port 456 nsew signal input
flabel metal2 s 192008 -800 192120 480 0 FreeSans 1120 90 0 0 la_oenb[18]
port 457 nsew signal input
flabel metal2 s 195554 -800 195666 480 0 FreeSans 1120 90 0 0 la_oenb[19]
port 458 nsew signal input
flabel metal2 s 131726 -800 131838 480 0 FreeSans 1120 90 0 0 la_oenb[1]
port 459 nsew signal input
flabel metal2 s 199100 -800 199212 480 0 FreeSans 1120 90 0 0 la_oenb[20]
port 460 nsew signal input
flabel metal2 s 202646 -800 202758 480 0 FreeSans 1120 90 0 0 la_oenb[21]
port 461 nsew signal input
flabel metal2 s 206192 -800 206304 480 0 FreeSans 1120 90 0 0 la_oenb[22]
port 462 nsew signal input
flabel metal2 s 209738 -800 209850 480 0 FreeSans 1120 90 0 0 la_oenb[23]
port 463 nsew signal input
flabel metal2 s 213284 -800 213396 480 0 FreeSans 1120 90 0 0 la_oenb[24]
port 464 nsew signal input
flabel metal2 s 216830 -800 216942 480 0 FreeSans 1120 90 0 0 la_oenb[25]
port 465 nsew signal input
flabel metal2 s 220376 -800 220488 480 0 FreeSans 1120 90 0 0 la_oenb[26]
port 466 nsew signal input
flabel metal2 s 223922 -800 224034 480 0 FreeSans 1120 90 0 0 la_oenb[27]
port 467 nsew signal input
flabel metal2 s 227468 -800 227580 480 0 FreeSans 1120 90 0 0 la_oenb[28]
port 468 nsew signal input
flabel metal2 s 231014 -800 231126 480 0 FreeSans 1120 90 0 0 la_oenb[29]
port 469 nsew signal input
flabel metal2 s 135272 -800 135384 480 0 FreeSans 1120 90 0 0 la_oenb[2]
port 470 nsew signal input
flabel metal2 s 234560 -800 234672 480 0 FreeSans 1120 90 0 0 la_oenb[30]
port 471 nsew signal input
flabel metal2 s 238106 -800 238218 480 0 FreeSans 1120 90 0 0 la_oenb[31]
port 472 nsew signal input
flabel metal2 s 241652 -800 241764 480 0 FreeSans 1120 90 0 0 la_oenb[32]
port 473 nsew signal input
flabel metal2 s 245198 -800 245310 480 0 FreeSans 1120 90 0 0 la_oenb[33]
port 474 nsew signal input
flabel metal2 s 248744 -800 248856 480 0 FreeSans 1120 90 0 0 la_oenb[34]
port 475 nsew signal input
flabel metal2 s 252290 -800 252402 480 0 FreeSans 1120 90 0 0 la_oenb[35]
port 476 nsew signal input
flabel metal2 s 255836 -800 255948 480 0 FreeSans 1120 90 0 0 la_oenb[36]
port 477 nsew signal input
flabel metal2 s 259382 -800 259494 480 0 FreeSans 1120 90 0 0 la_oenb[37]
port 478 nsew signal input
flabel metal2 s 262928 -800 263040 480 0 FreeSans 1120 90 0 0 la_oenb[38]
port 479 nsew signal input
flabel metal2 s 266474 -800 266586 480 0 FreeSans 1120 90 0 0 la_oenb[39]
port 480 nsew signal input
flabel metal2 s 138818 -800 138930 480 0 FreeSans 1120 90 0 0 la_oenb[3]
port 481 nsew signal input
flabel metal2 s 270020 -800 270132 480 0 FreeSans 1120 90 0 0 la_oenb[40]
port 482 nsew signal input
flabel metal2 s 273566 -800 273678 480 0 FreeSans 1120 90 0 0 la_oenb[41]
port 483 nsew signal input
flabel metal2 s 277112 -800 277224 480 0 FreeSans 1120 90 0 0 la_oenb[42]
port 484 nsew signal input
flabel metal2 s 280658 -800 280770 480 0 FreeSans 1120 90 0 0 la_oenb[43]
port 485 nsew signal input
flabel metal2 s 284204 -800 284316 480 0 FreeSans 1120 90 0 0 la_oenb[44]
port 486 nsew signal input
flabel metal2 s 287750 -800 287862 480 0 FreeSans 1120 90 0 0 la_oenb[45]
port 487 nsew signal input
flabel metal2 s 291296 -800 291408 480 0 FreeSans 1120 90 0 0 la_oenb[46]
port 488 nsew signal input
flabel metal2 s 294842 -800 294954 480 0 FreeSans 1120 90 0 0 la_oenb[47]
port 489 nsew signal input
flabel metal2 s 298388 -800 298500 480 0 FreeSans 1120 90 0 0 la_oenb[48]
port 490 nsew signal input
flabel metal2 s 301934 -800 302046 480 0 FreeSans 1120 90 0 0 la_oenb[49]
port 491 nsew signal input
flabel metal2 s 142364 -800 142476 480 0 FreeSans 1120 90 0 0 la_oenb[4]
port 492 nsew signal input
flabel metal2 s 305480 -800 305592 480 0 FreeSans 1120 90 0 0 la_oenb[50]
port 493 nsew signal input
flabel metal2 s 309026 -800 309138 480 0 FreeSans 1120 90 0 0 la_oenb[51]
port 494 nsew signal input
flabel metal2 s 312572 -800 312684 480 0 FreeSans 1120 90 0 0 la_oenb[52]
port 495 nsew signal input
flabel metal2 s 316118 -800 316230 480 0 FreeSans 1120 90 0 0 la_oenb[53]
port 496 nsew signal input
flabel metal2 s 319664 -800 319776 480 0 FreeSans 1120 90 0 0 la_oenb[54]
port 497 nsew signal input
flabel metal2 s 323210 -800 323322 480 0 FreeSans 1120 90 0 0 la_oenb[55]
port 498 nsew signal input
flabel metal2 s 326756 -800 326868 480 0 FreeSans 1120 90 0 0 la_oenb[56]
port 499 nsew signal input
flabel metal2 s 330302 -800 330414 480 0 FreeSans 1120 90 0 0 la_oenb[57]
port 500 nsew signal input
flabel metal2 s 333848 -800 333960 480 0 FreeSans 1120 90 0 0 la_oenb[58]
port 501 nsew signal input
flabel metal2 s 337394 -800 337506 480 0 FreeSans 1120 90 0 0 la_oenb[59]
port 502 nsew signal input
flabel metal2 s 145910 -800 146022 480 0 FreeSans 1120 90 0 0 la_oenb[5]
port 503 nsew signal input
flabel metal2 s 340940 -800 341052 480 0 FreeSans 1120 90 0 0 la_oenb[60]
port 504 nsew signal input
flabel metal2 s 344486 -800 344598 480 0 FreeSans 1120 90 0 0 la_oenb[61]
port 505 nsew signal input
flabel metal2 s 348032 -800 348144 480 0 FreeSans 1120 90 0 0 la_oenb[62]
port 506 nsew signal input
flabel metal2 s 351578 -800 351690 480 0 FreeSans 1120 90 0 0 la_oenb[63]
port 507 nsew signal input
flabel metal2 s 355124 -800 355236 480 0 FreeSans 1120 90 0 0 la_oenb[64]
port 508 nsew signal input
flabel metal2 s 358670 -800 358782 480 0 FreeSans 1120 90 0 0 la_oenb[65]
port 509 nsew signal input
flabel metal2 s 362216 -800 362328 480 0 FreeSans 1120 90 0 0 la_oenb[66]
port 510 nsew signal input
flabel metal2 s 365762 -800 365874 480 0 FreeSans 1120 90 0 0 la_oenb[67]
port 511 nsew signal input
flabel metal2 s 369308 -800 369420 480 0 FreeSans 1120 90 0 0 la_oenb[68]
port 512 nsew signal input
flabel metal2 s 372854 -800 372966 480 0 FreeSans 1120 90 0 0 la_oenb[69]
port 513 nsew signal input
flabel metal2 s 149456 -800 149568 480 0 FreeSans 1120 90 0 0 la_oenb[6]
port 514 nsew signal input
flabel metal2 s 376400 -800 376512 480 0 FreeSans 1120 90 0 0 la_oenb[70]
port 515 nsew signal input
flabel metal2 s 379946 -800 380058 480 0 FreeSans 1120 90 0 0 la_oenb[71]
port 516 nsew signal input
flabel metal2 s 383492 -800 383604 480 0 FreeSans 1120 90 0 0 la_oenb[72]
port 517 nsew signal input
flabel metal2 s 387038 -800 387150 480 0 FreeSans 1120 90 0 0 la_oenb[73]
port 518 nsew signal input
flabel metal2 s 390584 -800 390696 480 0 FreeSans 1120 90 0 0 la_oenb[74]
port 519 nsew signal input
flabel metal2 s 394130 -800 394242 480 0 FreeSans 1120 90 0 0 la_oenb[75]
port 520 nsew signal input
flabel metal2 s 397676 -800 397788 480 0 FreeSans 1120 90 0 0 la_oenb[76]
port 521 nsew signal input
flabel metal2 s 401222 -800 401334 480 0 FreeSans 1120 90 0 0 la_oenb[77]
port 522 nsew signal input
flabel metal2 s 404768 -800 404880 480 0 FreeSans 1120 90 0 0 la_oenb[78]
port 523 nsew signal input
flabel metal2 s 408314 -800 408426 480 0 FreeSans 1120 90 0 0 la_oenb[79]
port 524 nsew signal input
flabel metal2 s 153002 -800 153114 480 0 FreeSans 1120 90 0 0 la_oenb[7]
port 525 nsew signal input
flabel metal2 s 411860 -800 411972 480 0 FreeSans 1120 90 0 0 la_oenb[80]
port 526 nsew signal input
flabel metal2 s 415406 -800 415518 480 0 FreeSans 1120 90 0 0 la_oenb[81]
port 527 nsew signal input
flabel metal2 s 418952 -800 419064 480 0 FreeSans 1120 90 0 0 la_oenb[82]
port 528 nsew signal input
flabel metal2 s 422498 -800 422610 480 0 FreeSans 1120 90 0 0 la_oenb[83]
port 529 nsew signal input
flabel metal2 s 426044 -800 426156 480 0 FreeSans 1120 90 0 0 la_oenb[84]
port 530 nsew signal input
flabel metal2 s 429590 -800 429702 480 0 FreeSans 1120 90 0 0 la_oenb[85]
port 531 nsew signal input
flabel metal2 s 433136 -800 433248 480 0 FreeSans 1120 90 0 0 la_oenb[86]
port 532 nsew signal input
flabel metal2 s 436682 -800 436794 480 0 FreeSans 1120 90 0 0 la_oenb[87]
port 533 nsew signal input
flabel metal2 s 440228 -800 440340 480 0 FreeSans 1120 90 0 0 la_oenb[88]
port 534 nsew signal input
flabel metal2 s 443774 -800 443886 480 0 FreeSans 1120 90 0 0 la_oenb[89]
port 535 nsew signal input
flabel metal2 s 156548 -800 156660 480 0 FreeSans 1120 90 0 0 la_oenb[8]
port 536 nsew signal input
flabel metal2 s 447320 -800 447432 480 0 FreeSans 1120 90 0 0 la_oenb[90]
port 537 nsew signal input
flabel metal2 s 450866 -800 450978 480 0 FreeSans 1120 90 0 0 la_oenb[91]
port 538 nsew signal input
flabel metal2 s 454412 -800 454524 480 0 FreeSans 1120 90 0 0 la_oenb[92]
port 539 nsew signal input
flabel metal2 s 457958 -800 458070 480 0 FreeSans 1120 90 0 0 la_oenb[93]
port 540 nsew signal input
flabel metal2 s 461504 -800 461616 480 0 FreeSans 1120 90 0 0 la_oenb[94]
port 541 nsew signal input
flabel metal2 s 465050 -800 465162 480 0 FreeSans 1120 90 0 0 la_oenb[95]
port 542 nsew signal input
flabel metal2 s 468596 -800 468708 480 0 FreeSans 1120 90 0 0 la_oenb[96]
port 543 nsew signal input
flabel metal2 s 472142 -800 472254 480 0 FreeSans 1120 90 0 0 la_oenb[97]
port 544 nsew signal input
flabel metal2 s 475688 -800 475800 480 0 FreeSans 1120 90 0 0 la_oenb[98]
port 545 nsew signal input
flabel metal2 s 479234 -800 479346 480 0 FreeSans 1120 90 0 0 la_oenb[99]
port 546 nsew signal input
flabel metal2 s 160094 -800 160206 480 0 FreeSans 1120 90 0 0 la_oenb[9]
port 547 nsew signal input
flabel metal2 s 579704 -800 579816 480 0 FreeSans 1120 90 0 0 user_clock2
port 548 nsew signal input
flabel metal2 s 580886 -800 580998 480 0 FreeSans 1120 90 0 0 user_irq[0]
port 549 nsew signal tristate
flabel metal2 s 582068 -800 582180 480 0 FreeSans 1120 90 0 0 user_irq[1]
port 550 nsew signal tristate
flabel metal2 s 583250 -800 583362 480 0 FreeSans 1120 90 0 0 user_irq[2]
port 551 nsew signal tristate
flabel metal3 s 582340 639784 584800 644584 0 FreeSans 1120 0 0 0 vccd1
port 552 nsew signal bidirectional
flabel metal3 s 582340 629784 584800 634584 0 FreeSans 1120 0 0 0 vccd1
port 553 nsew signal bidirectional
flabel metal3 s 0 643842 1660 648642 0 FreeSans 1120 0 0 0 vccd2
port 554 nsew signal bidirectional
flabel metal3 s 0 633842 1660 638642 0 FreeSans 1120 0 0 0 vccd2
port 555 nsew signal bidirectional
flabel metal3 s 582340 540562 584800 545362 0 FreeSans 1120 0 0 0 vdda1
port 556 nsew signal bidirectional
flabel metal3 s 582340 550562 584800 555362 0 FreeSans 1120 0 0 0 vdda1
port 557 nsew signal bidirectional
flabel metal3 s 582340 235230 584800 240030 0 FreeSans 1120 0 0 0 vdda1
port 558 nsew signal bidirectional
flabel metal3 s 582340 225230 584800 230030 0 FreeSans 1120 0 0 0 vdda1
port 559 nsew signal bidirectional
flabel metal3 s 0 204888 1660 209688 0 FreeSans 1120 0 0 0 vdda2
port 560 nsew signal bidirectional
flabel metal3 s 0 214888 1660 219688 0 FreeSans 1120 0 0 0 vdda2
port 561 nsew signal bidirectional
flabel metal3 s 520594 702340 525394 704800 0 FreeSans 1920 180 0 0 vssa1
port 562 nsew signal bidirectional
flabel metal3 s 510594 702340 515394 704800 0 FreeSans 1920 180 0 0 vssa1
port 563 nsew signal bidirectional
flabel metal3 s 582340 146830 584800 151630 0 FreeSans 1120 0 0 0 vssa1
port 564 nsew signal bidirectional
flabel metal3 s 582340 136830 584800 141630 0 FreeSans 1120 0 0 0 vssa1
port 565 nsew signal bidirectional
flabel metal3 s 0 559442 1660 564242 0 FreeSans 1120 0 0 0 vssa2
port 566 nsew signal bidirectional
flabel metal3 s 0 549442 1660 554242 0 FreeSans 1120 0 0 0 vssa2
port 567 nsew signal bidirectional
flabel metal3 s 582340 191430 584800 196230 0 FreeSans 1120 0 0 0 vssd1
port 568 nsew signal bidirectional
flabel metal3 s 582340 181430 584800 186230 0 FreeSans 1120 0 0 0 vssd1
port 569 nsew signal bidirectional
flabel metal3 s 0 172888 1660 177688 0 FreeSans 1120 0 0 0 vssd2
port 570 nsew signal bidirectional
flabel metal3 s 0 162888 1660 167688 0 FreeSans 1120 0 0 0 vssd2
port 571 nsew signal bidirectional
flabel metal2 s 524 -800 636 480 0 FreeSans 1120 90 0 0 wb_clk_i
port 572 nsew signal input
flabel metal2 s 1706 -800 1818 480 0 FreeSans 1120 90 0 0 wb_rst_i
port 573 nsew signal input
flabel metal2 s 2888 -800 3000 480 0 FreeSans 1120 90 0 0 wbs_ack_o
port 574 nsew signal tristate
flabel metal2 s 7616 -800 7728 480 0 FreeSans 1120 90 0 0 wbs_adr_i[0]
port 575 nsew signal input
flabel metal2 s 47804 -800 47916 480 0 FreeSans 1120 90 0 0 wbs_adr_i[10]
port 576 nsew signal input
flabel metal2 s 51350 -800 51462 480 0 FreeSans 1120 90 0 0 wbs_adr_i[11]
port 577 nsew signal input
flabel metal2 s 54896 -800 55008 480 0 FreeSans 1120 90 0 0 wbs_adr_i[12]
port 578 nsew signal input
flabel metal2 s 58442 -800 58554 480 0 FreeSans 1120 90 0 0 wbs_adr_i[13]
port 579 nsew signal input
flabel metal2 s 61988 -800 62100 480 0 FreeSans 1120 90 0 0 wbs_adr_i[14]
port 580 nsew signal input
flabel metal2 s 65534 -800 65646 480 0 FreeSans 1120 90 0 0 wbs_adr_i[15]
port 581 nsew signal input
flabel metal2 s 69080 -800 69192 480 0 FreeSans 1120 90 0 0 wbs_adr_i[16]
port 582 nsew signal input
flabel metal2 s 72626 -800 72738 480 0 FreeSans 1120 90 0 0 wbs_adr_i[17]
port 583 nsew signal input
flabel metal2 s 76172 -800 76284 480 0 FreeSans 1120 90 0 0 wbs_adr_i[18]
port 584 nsew signal input
flabel metal2 s 79718 -800 79830 480 0 FreeSans 1120 90 0 0 wbs_adr_i[19]
port 585 nsew signal input
flabel metal2 s 12344 -800 12456 480 0 FreeSans 1120 90 0 0 wbs_adr_i[1]
port 586 nsew signal input
flabel metal2 s 83264 -800 83376 480 0 FreeSans 1120 90 0 0 wbs_adr_i[20]
port 587 nsew signal input
flabel metal2 s 86810 -800 86922 480 0 FreeSans 1120 90 0 0 wbs_adr_i[21]
port 588 nsew signal input
flabel metal2 s 90356 -800 90468 480 0 FreeSans 1120 90 0 0 wbs_adr_i[22]
port 589 nsew signal input
flabel metal2 s 93902 -800 94014 480 0 FreeSans 1120 90 0 0 wbs_adr_i[23]
port 590 nsew signal input
flabel metal2 s 97448 -800 97560 480 0 FreeSans 1120 90 0 0 wbs_adr_i[24]
port 591 nsew signal input
flabel metal2 s 100994 -800 101106 480 0 FreeSans 1120 90 0 0 wbs_adr_i[25]
port 592 nsew signal input
flabel metal2 s 104540 -800 104652 480 0 FreeSans 1120 90 0 0 wbs_adr_i[26]
port 593 nsew signal input
flabel metal2 s 108086 -800 108198 480 0 FreeSans 1120 90 0 0 wbs_adr_i[27]
port 594 nsew signal input
flabel metal2 s 111632 -800 111744 480 0 FreeSans 1120 90 0 0 wbs_adr_i[28]
port 595 nsew signal input
flabel metal2 s 115178 -800 115290 480 0 FreeSans 1120 90 0 0 wbs_adr_i[29]
port 596 nsew signal input
flabel metal2 s 17072 -800 17184 480 0 FreeSans 1120 90 0 0 wbs_adr_i[2]
port 597 nsew signal input
flabel metal2 s 118724 -800 118836 480 0 FreeSans 1120 90 0 0 wbs_adr_i[30]
port 598 nsew signal input
flabel metal2 s 122270 -800 122382 480 0 FreeSans 1120 90 0 0 wbs_adr_i[31]
port 599 nsew signal input
flabel metal2 s 21800 -800 21912 480 0 FreeSans 1120 90 0 0 wbs_adr_i[3]
port 600 nsew signal input
flabel metal2 s 26528 -800 26640 480 0 FreeSans 1120 90 0 0 wbs_adr_i[4]
port 601 nsew signal input
flabel metal2 s 30074 -800 30186 480 0 FreeSans 1120 90 0 0 wbs_adr_i[5]
port 602 nsew signal input
flabel metal2 s 33620 -800 33732 480 0 FreeSans 1120 90 0 0 wbs_adr_i[6]
port 603 nsew signal input
flabel metal2 s 37166 -800 37278 480 0 FreeSans 1120 90 0 0 wbs_adr_i[7]
port 604 nsew signal input
flabel metal2 s 40712 -800 40824 480 0 FreeSans 1120 90 0 0 wbs_adr_i[8]
port 605 nsew signal input
flabel metal2 s 44258 -800 44370 480 0 FreeSans 1120 90 0 0 wbs_adr_i[9]
port 606 nsew signal input
flabel metal2 s 4070 -800 4182 480 0 FreeSans 1120 90 0 0 wbs_cyc_i
port 607 nsew signal input
flabel metal2 s 8798 -800 8910 480 0 FreeSans 1120 90 0 0 wbs_dat_i[0]
port 608 nsew signal input
flabel metal2 s 48986 -800 49098 480 0 FreeSans 1120 90 0 0 wbs_dat_i[10]
port 609 nsew signal input
flabel metal2 s 52532 -800 52644 480 0 FreeSans 1120 90 0 0 wbs_dat_i[11]
port 610 nsew signal input
flabel metal2 s 56078 -800 56190 480 0 FreeSans 1120 90 0 0 wbs_dat_i[12]
port 611 nsew signal input
flabel metal2 s 59624 -800 59736 480 0 FreeSans 1120 90 0 0 wbs_dat_i[13]
port 612 nsew signal input
flabel metal2 s 63170 -800 63282 480 0 FreeSans 1120 90 0 0 wbs_dat_i[14]
port 613 nsew signal input
flabel metal2 s 66716 -800 66828 480 0 FreeSans 1120 90 0 0 wbs_dat_i[15]
port 614 nsew signal input
flabel metal2 s 70262 -800 70374 480 0 FreeSans 1120 90 0 0 wbs_dat_i[16]
port 615 nsew signal input
flabel metal2 s 73808 -800 73920 480 0 FreeSans 1120 90 0 0 wbs_dat_i[17]
port 616 nsew signal input
flabel metal2 s 77354 -800 77466 480 0 FreeSans 1120 90 0 0 wbs_dat_i[18]
port 617 nsew signal input
flabel metal2 s 80900 -800 81012 480 0 FreeSans 1120 90 0 0 wbs_dat_i[19]
port 618 nsew signal input
flabel metal2 s 13526 -800 13638 480 0 FreeSans 1120 90 0 0 wbs_dat_i[1]
port 619 nsew signal input
flabel metal2 s 84446 -800 84558 480 0 FreeSans 1120 90 0 0 wbs_dat_i[20]
port 620 nsew signal input
flabel metal2 s 87992 -800 88104 480 0 FreeSans 1120 90 0 0 wbs_dat_i[21]
port 621 nsew signal input
flabel metal2 s 91538 -800 91650 480 0 FreeSans 1120 90 0 0 wbs_dat_i[22]
port 622 nsew signal input
flabel metal2 s 95084 -800 95196 480 0 FreeSans 1120 90 0 0 wbs_dat_i[23]
port 623 nsew signal input
flabel metal2 s 98630 -800 98742 480 0 FreeSans 1120 90 0 0 wbs_dat_i[24]
port 624 nsew signal input
flabel metal2 s 102176 -800 102288 480 0 FreeSans 1120 90 0 0 wbs_dat_i[25]
port 625 nsew signal input
flabel metal2 s 105722 -800 105834 480 0 FreeSans 1120 90 0 0 wbs_dat_i[26]
port 626 nsew signal input
flabel metal2 s 109268 -800 109380 480 0 FreeSans 1120 90 0 0 wbs_dat_i[27]
port 627 nsew signal input
flabel metal2 s 112814 -800 112926 480 0 FreeSans 1120 90 0 0 wbs_dat_i[28]
port 628 nsew signal input
flabel metal2 s 116360 -800 116472 480 0 FreeSans 1120 90 0 0 wbs_dat_i[29]
port 629 nsew signal input
flabel metal2 s 18254 -800 18366 480 0 FreeSans 1120 90 0 0 wbs_dat_i[2]
port 630 nsew signal input
flabel metal2 s 119906 -800 120018 480 0 FreeSans 1120 90 0 0 wbs_dat_i[30]
port 631 nsew signal input
flabel metal2 s 123452 -800 123564 480 0 FreeSans 1120 90 0 0 wbs_dat_i[31]
port 632 nsew signal input
flabel metal2 s 22982 -800 23094 480 0 FreeSans 1120 90 0 0 wbs_dat_i[3]
port 633 nsew signal input
flabel metal2 s 27710 -800 27822 480 0 FreeSans 1120 90 0 0 wbs_dat_i[4]
port 634 nsew signal input
flabel metal2 s 31256 -800 31368 480 0 FreeSans 1120 90 0 0 wbs_dat_i[5]
port 635 nsew signal input
flabel metal2 s 34802 -800 34914 480 0 FreeSans 1120 90 0 0 wbs_dat_i[6]
port 636 nsew signal input
flabel metal2 s 38348 -800 38460 480 0 FreeSans 1120 90 0 0 wbs_dat_i[7]
port 637 nsew signal input
flabel metal2 s 41894 -800 42006 480 0 FreeSans 1120 90 0 0 wbs_dat_i[8]
port 638 nsew signal input
flabel metal2 s 45440 -800 45552 480 0 FreeSans 1120 90 0 0 wbs_dat_i[9]
port 639 nsew signal input
flabel metal2 s 9980 -800 10092 480 0 FreeSans 1120 90 0 0 wbs_dat_o[0]
port 640 nsew signal tristate
flabel metal2 s 50168 -800 50280 480 0 FreeSans 1120 90 0 0 wbs_dat_o[10]
port 641 nsew signal tristate
flabel metal2 s 53714 -800 53826 480 0 FreeSans 1120 90 0 0 wbs_dat_o[11]
port 642 nsew signal tristate
flabel metal2 s 57260 -800 57372 480 0 FreeSans 1120 90 0 0 wbs_dat_o[12]
port 643 nsew signal tristate
flabel metal2 s 60806 -800 60918 480 0 FreeSans 1120 90 0 0 wbs_dat_o[13]
port 644 nsew signal tristate
flabel metal2 s 64352 -800 64464 480 0 FreeSans 1120 90 0 0 wbs_dat_o[14]
port 645 nsew signal tristate
flabel metal2 s 67898 -800 68010 480 0 FreeSans 1120 90 0 0 wbs_dat_o[15]
port 646 nsew signal tristate
flabel metal2 s 71444 -800 71556 480 0 FreeSans 1120 90 0 0 wbs_dat_o[16]
port 647 nsew signal tristate
flabel metal2 s 74990 -800 75102 480 0 FreeSans 1120 90 0 0 wbs_dat_o[17]
port 648 nsew signal tristate
flabel metal2 s 78536 -800 78648 480 0 FreeSans 1120 90 0 0 wbs_dat_o[18]
port 649 nsew signal tristate
flabel metal2 s 82082 -800 82194 480 0 FreeSans 1120 90 0 0 wbs_dat_o[19]
port 650 nsew signal tristate
flabel metal2 s 14708 -800 14820 480 0 FreeSans 1120 90 0 0 wbs_dat_o[1]
port 651 nsew signal tristate
flabel metal2 s 85628 -800 85740 480 0 FreeSans 1120 90 0 0 wbs_dat_o[20]
port 652 nsew signal tristate
flabel metal2 s 89174 -800 89286 480 0 FreeSans 1120 90 0 0 wbs_dat_o[21]
port 653 nsew signal tristate
flabel metal2 s 92720 -800 92832 480 0 FreeSans 1120 90 0 0 wbs_dat_o[22]
port 654 nsew signal tristate
flabel metal2 s 96266 -800 96378 480 0 FreeSans 1120 90 0 0 wbs_dat_o[23]
port 655 nsew signal tristate
flabel metal2 s 99812 -800 99924 480 0 FreeSans 1120 90 0 0 wbs_dat_o[24]
port 656 nsew signal tristate
flabel metal2 s 103358 -800 103470 480 0 FreeSans 1120 90 0 0 wbs_dat_o[25]
port 657 nsew signal tristate
flabel metal2 s 106904 -800 107016 480 0 FreeSans 1120 90 0 0 wbs_dat_o[26]
port 658 nsew signal tristate
flabel metal2 s 110450 -800 110562 480 0 FreeSans 1120 90 0 0 wbs_dat_o[27]
port 659 nsew signal tristate
flabel metal2 s 113996 -800 114108 480 0 FreeSans 1120 90 0 0 wbs_dat_o[28]
port 660 nsew signal tristate
flabel metal2 s 117542 -800 117654 480 0 FreeSans 1120 90 0 0 wbs_dat_o[29]
port 661 nsew signal tristate
flabel metal2 s 19436 -800 19548 480 0 FreeSans 1120 90 0 0 wbs_dat_o[2]
port 662 nsew signal tristate
flabel metal2 s 121088 -800 121200 480 0 FreeSans 1120 90 0 0 wbs_dat_o[30]
port 663 nsew signal tristate
flabel metal2 s 124634 -800 124746 480 0 FreeSans 1120 90 0 0 wbs_dat_o[31]
port 664 nsew signal tristate
flabel metal2 s 24164 -800 24276 480 0 FreeSans 1120 90 0 0 wbs_dat_o[3]
port 665 nsew signal tristate
flabel metal2 s 28892 -800 29004 480 0 FreeSans 1120 90 0 0 wbs_dat_o[4]
port 666 nsew signal tristate
flabel metal2 s 32438 -800 32550 480 0 FreeSans 1120 90 0 0 wbs_dat_o[5]
port 667 nsew signal tristate
flabel metal2 s 35984 -800 36096 480 0 FreeSans 1120 90 0 0 wbs_dat_o[6]
port 668 nsew signal tristate
flabel metal2 s 39530 -800 39642 480 0 FreeSans 1120 90 0 0 wbs_dat_o[7]
port 669 nsew signal tristate
flabel metal2 s 43076 -800 43188 480 0 FreeSans 1120 90 0 0 wbs_dat_o[8]
port 670 nsew signal tristate
flabel metal2 s 46622 -800 46734 480 0 FreeSans 1120 90 0 0 wbs_dat_o[9]
port 671 nsew signal tristate
flabel metal2 s 11162 -800 11274 480 0 FreeSans 1120 90 0 0 wbs_sel_i[0]
port 672 nsew signal input
flabel metal2 s 15890 -800 16002 480 0 FreeSans 1120 90 0 0 wbs_sel_i[1]
port 673 nsew signal input
flabel metal2 s 20618 -800 20730 480 0 FreeSans 1120 90 0 0 wbs_sel_i[2]
port 674 nsew signal input
flabel metal2 s 25346 -800 25458 480 0 FreeSans 1120 90 0 0 wbs_sel_i[3]
port 675 nsew signal input
flabel metal2 s 5252 -800 5364 480 0 FreeSans 1120 90 0 0 wbs_stb_i
port 676 nsew signal input
flabel metal2 s 6434 -800 6546 480 0 FreeSans 1120 90 0 0 wbs_we_i
port 677 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
